module alu (carry_out,
    clk,
    overflow,
    zero,
    alu_op,
    op1,
    op2,
    result);
 output carry_out;
 input clk;
 output overflow;
 output zero;
 input [3:0] alu_op;
 input [31:0] op1;
 input [31:0] op2;
 output [31:0] result;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire net103;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;

 sky130_fd_sc_hd__clkbuf_4 _0982_ (.A(net63),
    .X(_0018_));
 sky130_fd_sc_hd__clkbuf_4 _0983_ (.A(net37),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _0984_ (.A0(net25),
    .A1(net26),
    .S(_0029_),
    .X(_0039_));
 sky130_fd_sc_hd__buf_2 _0985_ (.A(net28),
    .X(_0050_));
 sky130_fd_sc_hd__buf_2 _0986_ (.A(net29),
    .X(_0060_));
 sky130_fd_sc_hd__buf_4 _0987_ (.A(_0029_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _0988_ (.A0(_0050_),
    .A1(_0060_),
    .S(_0071_),
    .X(_0081_));
 sky130_fd_sc_hd__clkbuf_4 _0989_ (.A(net48),
    .X(_0091_));
 sky130_fd_sc_hd__clkbuf_4 _0990_ (.A(_0091_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _0991_ (.A0(_0039_),
    .A1(_0081_),
    .S(_0102_),
    .X(_0112_));
 sky130_fd_sc_hd__buf_2 _0992_ (.A(net23),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _0993_ (.A0(_0119_),
    .A1(net24),
    .S(_0029_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _0994_ (.A0(net21),
    .A1(net22),
    .S(_0029_),
    .X(_0121_));
 sky130_fd_sc_hd__inv_2 _0995_ (.A(_0091_),
    .Y(_0122_));
 sky130_fd_sc_hd__mux2_1 _0996_ (.A0(_0120_),
    .A1(_0121_),
    .S(_0122_),
    .X(_0123_));
 sky130_fd_sc_hd__clkbuf_4 _0997_ (.A(net59),
    .X(_0124_));
 sky130_fd_sc_hd__inv_2 _0998_ (.A(_0124_),
    .Y(_0125_));
 sky130_fd_sc_hd__clkbuf_4 _0999_ (.A(_0125_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _1000_ (.A0(_0112_),
    .A1(_0123_),
    .S(_0126_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _1001_ (.A0(net19),
    .A1(net20),
    .S(_0029_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _1002_ (.A0(net17),
    .A1(net18),
    .S(_0029_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _1003_ (.A0(_0128_),
    .A1(_0129_),
    .S(_0122_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _1004_ (.A0(net14),
    .A1(net15),
    .S(_0071_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _1005_ (.A0(net12),
    .A1(net13),
    .S(_0071_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _1006_ (.A0(_0131_),
    .A1(_0132_),
    .S(_0122_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _1007_ (.A0(_0130_),
    .A1(_0133_),
    .S(_0125_),
    .X(_0134_));
 sky130_fd_sc_hd__clkbuf_4 _1008_ (.A(net62),
    .X(_0135_));
 sky130_fd_sc_hd__inv_2 _1009_ (.A(_0135_),
    .Y(_0136_));
 sky130_fd_sc_hd__buf_2 _1010_ (.A(_0136_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _1011_ (.A0(_0127_),
    .A1(_0134_),
    .S(_0137_),
    .X(_0138_));
 sky130_fd_sc_hd__clkbuf_2 _1012_ (.A(net4),
    .X(_0139_));
 sky130_fd_sc_hd__clkbuf_2 _1013_ (.A(net3),
    .X(_0140_));
 sky130_fd_sc_hd__buf_2 _1014_ (.A(net2),
    .X(_0141_));
 sky130_fd_sc_hd__and3b_2 _1015_ (.A_N(_0139_),
    .B(_0140_),
    .C(_0141_),
    .X(_0142_));
 sky130_fd_sc_hd__buf_2 _1016_ (.A(net9),
    .X(_0143_));
 sky130_fd_sc_hd__buf_4 _1017_ (.A(_0029_),
    .X(_0144_));
 sky130_fd_sc_hd__mux4_1 _1018_ (.A0(net8),
    .A1(_0143_),
    .A2(net10),
    .A3(net11),
    .S0(_0144_),
    .S1(_0091_),
    .X(_0145_));
 sky130_fd_sc_hd__clkbuf_2 _1019_ (.A(net36),
    .X(_0146_));
 sky130_fd_sc_hd__clkbuf_2 _1020_ (.A(net7),
    .X(_0147_));
 sky130_fd_sc_hd__mux4_1 _1021_ (.A0(net35),
    .A1(_0146_),
    .A2(net6),
    .A3(_0147_),
    .S0(_0144_),
    .S1(_0091_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _1022_ (.A0(_0145_),
    .A1(_0148_),
    .S(_0125_),
    .X(_0149_));
 sky130_fd_sc_hd__nor2_2 _1023_ (.A(net48),
    .B(net37),
    .Y(_0150_));
 sky130_fd_sc_hd__nand2_2 _1024_ (.A(net5),
    .B(_0150_),
    .Y(_0151_));
 sky130_fd_sc_hd__nor2_2 _1025_ (.A(_0135_),
    .B(_0124_),
    .Y(_0152_));
 sky130_fd_sc_hd__nand2_1 _1026_ (.A(_0151_),
    .B(_0152_),
    .Y(_0153_));
 sky130_fd_sc_hd__buf_2 _1027_ (.A(_0102_),
    .X(_0154_));
 sky130_fd_sc_hd__buf_2 _1028_ (.A(net27),
    .X(_0155_));
 sky130_fd_sc_hd__buf_2 _1029_ (.A(net30),
    .X(_0156_));
 sky130_fd_sc_hd__clkbuf_4 _1030_ (.A(_0071_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _1031_ (.A0(_0155_),
    .A1(_0156_),
    .S(_0157_),
    .X(_0158_));
 sky130_fd_sc_hd__buf_2 _1032_ (.A(net16),
    .X(_0159_));
 sky130_fd_sc_hd__clkbuf_4 _1033_ (.A(_0122_),
    .X(_0160_));
 sky130_fd_sc_hd__and3_1 _1034_ (.A(_0159_),
    .B(_0160_),
    .C(_0157_),
    .X(_0161_));
 sky130_fd_sc_hd__a21o_1 _1035_ (.A1(_0154_),
    .A2(_0158_),
    .B1(_0161_),
    .X(_0162_));
 sky130_fd_sc_hd__nand2_1 _1036_ (.A(_0136_),
    .B(_0124_),
    .Y(_0163_));
 sky130_fd_sc_hd__buf_2 _1037_ (.A(net31),
    .X(_0164_));
 sky130_fd_sc_hd__clkbuf_2 _1038_ (.A(net32),
    .X(_0165_));
 sky130_fd_sc_hd__clkbuf_2 _1039_ (.A(net33),
    .X(_0166_));
 sky130_fd_sc_hd__buf_2 _1040_ (.A(net34),
    .X(_0167_));
 sky130_fd_sc_hd__mux4_1 _1041_ (.A0(_0164_),
    .A1(_0165_),
    .A2(_0166_),
    .A3(_0167_),
    .S0(_0157_),
    .S1(_0102_),
    .X(_0168_));
 sky130_fd_sc_hd__o22a_1 _1042_ (.A1(_0153_),
    .A2(_0162_),
    .B1(_0163_),
    .B2(_0168_),
    .X(_0169_));
 sky130_fd_sc_hd__nand3b_2 _1043_ (.A_N(_0139_),
    .B(_0140_),
    .C(net2),
    .Y(_0170_));
 sky130_fd_sc_hd__nor2_2 _1044_ (.A(_0018_),
    .B(_0170_),
    .Y(_0171_));
 sky130_fd_sc_hd__o211a_1 _1045_ (.A1(_0137_),
    .A2(_0149_),
    .B1(_0169_),
    .C1(_0171_),
    .X(_0172_));
 sky130_fd_sc_hd__or4bb_2 _1046_ (.A(net2),
    .B(_0139_),
    .C_N(_0140_),
    .D_N(net1),
    .X(_0173_));
 sky130_fd_sc_hd__nor2_2 _1047_ (.A(_0018_),
    .B(_0173_),
    .Y(_0174_));
 sky130_fd_sc_hd__nand2_1 _1048_ (.A(_0174_),
    .B(_0152_),
    .Y(_0175_));
 sky130_fd_sc_hd__buf_4 _1049_ (.A(_0071_),
    .X(_0176_));
 sky130_fd_sc_hd__nor2_1 _1050_ (.A(net5),
    .B(_0176_),
    .Y(_0177_));
 sky130_fd_sc_hd__nor2_2 _1051_ (.A(_0140_),
    .B(_0139_),
    .Y(_0178_));
 sky130_fd_sc_hd__nand3_4 _1052_ (.A(net1),
    .B(_0141_),
    .C(_0178_),
    .Y(_0179_));
 sky130_fd_sc_hd__and2_1 _1053_ (.A(net5),
    .B(_0071_),
    .X(_0180_));
 sky130_fd_sc_hd__inv_2 _1054_ (.A(net1),
    .Y(_0181_));
 sky130_fd_sc_hd__and3_1 _1055_ (.A(_0181_),
    .B(net2),
    .C(_0178_),
    .X(_0182_));
 sky130_fd_sc_hd__nand2_1 _1056_ (.A(_0180_),
    .B(_0182_),
    .Y(_0183_));
 sky130_fd_sc_hd__or3_1 _1057_ (.A(net2),
    .B(_0140_),
    .C(_0139_),
    .X(_0184_));
 sky130_fd_sc_hd__clkbuf_4 _1058_ (.A(_0184_),
    .X(_0185_));
 sky130_fd_sc_hd__or4b_1 _1059_ (.A(net1),
    .B(net2),
    .C(_0139_),
    .D_N(_0140_),
    .X(_0186_));
 sky130_fd_sc_hd__a211o_1 _1060_ (.A1(_0185_),
    .A2(_0186_),
    .B1(_0180_),
    .C1(_0177_),
    .X(_0187_));
 sky130_fd_sc_hd__o211a_1 _1061_ (.A1(_0177_),
    .A2(_0179_),
    .B1(_0183_),
    .C1(_0187_),
    .X(_0188_));
 sky130_fd_sc_hd__o21a_1 _1062_ (.A1(_0151_),
    .A2(_0175_),
    .B1(_0188_),
    .X(_0189_));
 sky130_fd_sc_hd__inv_2 _1063_ (.A(_0189_),
    .Y(_0190_));
 sky130_fd_sc_hd__a311o_1 _1064_ (.A1(_0018_),
    .A2(_0138_),
    .A3(_0142_),
    .B1(_0172_),
    .C1(_0190_),
    .X(_0191_));
 sky130_fd_sc_hd__inv_2 _1065_ (.A(net5),
    .Y(_0192_));
 sky130_fd_sc_hd__clkbuf_4 _1066_ (.A(_0091_),
    .X(_0193_));
 sky130_fd_sc_hd__o21ai_1 _1067_ (.A1(_0192_),
    .A2(_0176_),
    .B1(_0193_),
    .Y(_0194_));
 sky130_fd_sc_hd__or2_1 _1068_ (.A(net30),
    .B(net62),
    .X(_0195_));
 sky130_fd_sc_hd__nand2_1 _1069_ (.A(net30),
    .B(_0135_),
    .Y(_0196_));
 sky130_fd_sc_hd__or2_1 _1070_ (.A(net27),
    .B(net59),
    .X(_0197_));
 sky130_fd_sc_hd__nand2_1 _1071_ (.A(net27),
    .B(_0124_),
    .Y(_0198_));
 sky130_fd_sc_hd__a22o_1 _1072_ (.A1(_0195_),
    .A2(_0196_),
    .B1(_0197_),
    .B2(_0198_),
    .X(_0199_));
 sky130_fd_sc_hd__a221o_1 _1073_ (.A1(net5),
    .A2(_0150_),
    .B1(_0194_),
    .B2(_0159_),
    .C1(_0199_),
    .X(_0200_));
 sky130_fd_sc_hd__a211o_1 _1074_ (.A1(_0195_),
    .A2(_0196_),
    .B1(_0155_),
    .C1(_0125_),
    .X(_0201_));
 sky130_fd_sc_hd__or2_1 _1075_ (.A(_0156_),
    .B(_0136_),
    .X(_0202_));
 sky130_fd_sc_hd__nand2_1 _1076_ (.A(net33),
    .B(net65),
    .Y(_0203_));
 sky130_fd_sc_hd__or2_1 _1077_ (.A(net33),
    .B(net65),
    .X(_0204_));
 sky130_fd_sc_hd__xor2_2 _1078_ (.A(net34),
    .B(net66),
    .X(_0205_));
 sky130_fd_sc_hd__a21oi_1 _1079_ (.A1(_0203_),
    .A2(_0204_),
    .B1(_0205_),
    .Y(_0206_));
 sky130_fd_sc_hd__nand2_1 _1080_ (.A(net32),
    .B(net64),
    .Y(_0207_));
 sky130_fd_sc_hd__or2_1 _1081_ (.A(net32),
    .B(net64),
    .X(_0208_));
 sky130_fd_sc_hd__nand2_1 _1082_ (.A(_0207_),
    .B(_0208_),
    .Y(_0209_));
 sky130_fd_sc_hd__nand2_1 _1083_ (.A(_0018_),
    .B(_0164_),
    .Y(_0210_));
 sky130_fd_sc_hd__or2_1 _1084_ (.A(_0018_),
    .B(net31),
    .X(_0211_));
 sky130_fd_sc_hd__nand2_1 _1085_ (.A(_0210_),
    .B(_0211_),
    .Y(_0212_));
 sky130_fd_sc_hd__nand3_1 _1086_ (.A(_0206_),
    .B(_0209_),
    .C(_0212_),
    .Y(_0213_));
 sky130_fd_sc_hd__a31o_1 _1087_ (.A1(_0200_),
    .A2(_0201_),
    .A3(_0202_),
    .B1(_0213_),
    .X(_0214_));
 sky130_fd_sc_hd__or3b_1 _1088_ (.A(_0166_),
    .B(_0205_),
    .C_N(net65),
    .X(_0215_));
 sky130_fd_sc_hd__inv_2 _1089_ (.A(_0164_),
    .Y(_0216_));
 sky130_fd_sc_hd__inv_2 _1090_ (.A(net32),
    .Y(_0217_));
 sky130_fd_sc_hd__and2_1 _1091_ (.A(_0217_),
    .B(net64),
    .X(_0218_));
 sky130_fd_sc_hd__a31o_1 _1092_ (.A1(_0018_),
    .A2(_0216_),
    .A3(_0209_),
    .B1(_0218_),
    .X(_0219_));
 sky130_fd_sc_hd__inv_2 _1093_ (.A(net66),
    .Y(_0220_));
 sky130_fd_sc_hd__o2bb2a_1 _1094_ (.A1_N(_0206_),
    .A2_N(_0219_),
    .B1(_0167_),
    .B2(_0220_),
    .X(_0221_));
 sky130_fd_sc_hd__xor2_1 _1095_ (.A(net9),
    .B(net41),
    .X(_0222_));
 sky130_fd_sc_hd__or2_1 _1096_ (.A(net40),
    .B(net8),
    .X(_0223_));
 sky130_fd_sc_hd__nand2_1 _1097_ (.A(net40),
    .B(net8),
    .Y(_0224_));
 sky130_fd_sc_hd__and2_1 _1098_ (.A(_0223_),
    .B(_0224_),
    .X(_0225_));
 sky130_fd_sc_hd__xnor2_1 _1099_ (.A(net11),
    .B(net43),
    .Y(_0226_));
 sky130_fd_sc_hd__xnor2_1 _1100_ (.A(net10),
    .B(net42),
    .Y(_0227_));
 sky130_fd_sc_hd__and2_1 _1101_ (.A(_0226_),
    .B(_0227_),
    .X(_0228_));
 sky130_fd_sc_hd__or3b_1 _1102_ (.A(_0222_),
    .B(_0225_),
    .C_N(_0228_),
    .X(_0229_));
 sky130_fd_sc_hd__xor2_1 _1103_ (.A(net36),
    .B(net68),
    .X(_0230_));
 sky130_fd_sc_hd__and2_1 _1104_ (.A(net67),
    .B(net35),
    .X(_0231_));
 sky130_fd_sc_hd__clkbuf_2 _1105_ (.A(net35),
    .X(_0232_));
 sky130_fd_sc_hd__nor2_1 _1106_ (.A(net67),
    .B(_0232_),
    .Y(_0233_));
 sky130_fd_sc_hd__nor2_1 _1107_ (.A(_0231_),
    .B(_0233_),
    .Y(_0234_));
 sky130_fd_sc_hd__or2_1 _1108_ (.A(net6),
    .B(net38),
    .X(_0235_));
 sky130_fd_sc_hd__nand2_1 _1109_ (.A(net6),
    .B(net38),
    .Y(_0236_));
 sky130_fd_sc_hd__nor2_1 _1110_ (.A(net7),
    .B(net39),
    .Y(_0237_));
 sky130_fd_sc_hd__and2_1 _1111_ (.A(net7),
    .B(net39),
    .X(_0238_));
 sky130_fd_sc_hd__nor2_1 _1112_ (.A(_0237_),
    .B(_0238_),
    .Y(_0239_));
 sky130_fd_sc_hd__a21oi_1 _1113_ (.A1(_0235_),
    .A2(_0236_),
    .B1(_0239_),
    .Y(_0240_));
 sky130_fd_sc_hd__or4b_2 _1114_ (.A(_0229_),
    .B(_0230_),
    .C(_0234_),
    .D_N(_0240_),
    .X(_0241_));
 sky130_fd_sc_hd__a31o_1 _1115_ (.A1(_0214_),
    .A2(_0215_),
    .A3(_0221_),
    .B1(_0241_),
    .X(_0242_));
 sky130_fd_sc_hd__buf_2 _1116_ (.A(net11),
    .X(_0243_));
 sky130_fd_sc_hd__inv_2 _1117_ (.A(net43),
    .Y(_0244_));
 sky130_fd_sc_hd__buf_2 _1118_ (.A(net10),
    .X(_0245_));
 sky130_fd_sc_hd__nand2_1 _1119_ (.A(net42),
    .B(_0226_),
    .Y(_0246_));
 sky130_fd_sc_hd__inv_2 _1120_ (.A(_0143_),
    .Y(_0247_));
 sky130_fd_sc_hd__clkbuf_2 _1121_ (.A(net8),
    .X(_0248_));
 sky130_fd_sc_hd__nor2_1 _1122_ (.A(_0248_),
    .B(_0222_),
    .Y(_0249_));
 sky130_fd_sc_hd__a22o_1 _1123_ (.A1(_0247_),
    .A2(net41),
    .B1(net40),
    .B2(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__nand2_1 _1124_ (.A(_0228_),
    .B(_0250_),
    .Y(_0251_));
 sky130_fd_sc_hd__o221a_1 _1125_ (.A1(_0243_),
    .A2(_0244_),
    .B1(_0245_),
    .B2(_0246_),
    .C1(_0251_),
    .X(_0252_));
 sky130_fd_sc_hd__clkbuf_2 _1126_ (.A(net6),
    .X(_0253_));
 sky130_fd_sc_hd__or3b_1 _1127_ (.A(_0253_),
    .B(_0239_),
    .C_N(net38),
    .X(_0254_));
 sky130_fd_sc_hd__inv_2 _1128_ (.A(net36),
    .Y(_0255_));
 sky130_fd_sc_hd__nor2_1 _1129_ (.A(_0232_),
    .B(_0230_),
    .Y(_0256_));
 sky130_fd_sc_hd__a22o_1 _1130_ (.A1(_0255_),
    .A2(net68),
    .B1(net67),
    .B2(_0256_),
    .X(_0257_));
 sky130_fd_sc_hd__inv_2 _1131_ (.A(net39),
    .Y(_0258_));
 sky130_fd_sc_hd__o2bb2a_1 _1132_ (.A1_N(_0240_),
    .A2_N(_0257_),
    .B1(_0147_),
    .B2(_0258_),
    .X(_0259_));
 sky130_fd_sc_hd__a21o_1 _1133_ (.A1(_0254_),
    .A2(_0259_),
    .B1(_0229_),
    .X(_0260_));
 sky130_fd_sc_hd__or2_1 _1134_ (.A(net53),
    .B(net21),
    .X(_0261_));
 sky130_fd_sc_hd__nand2_1 _1135_ (.A(net53),
    .B(net21),
    .Y(_0262_));
 sky130_fd_sc_hd__and2_1 _1136_ (.A(_0261_),
    .B(_0262_),
    .X(_0263_));
 sky130_fd_sc_hd__or2_1 _1137_ (.A(net24),
    .B(net56),
    .X(_0264_));
 sky130_fd_sc_hd__nand2_1 _1138_ (.A(net24),
    .B(net56),
    .Y(_0265_));
 sky130_fd_sc_hd__or2_1 _1139_ (.A(net23),
    .B(net55),
    .X(_0266_));
 sky130_fd_sc_hd__nand2_1 _1140_ (.A(net23),
    .B(net55),
    .Y(_0267_));
 sky130_fd_sc_hd__a22o_1 _1141_ (.A1(_0264_),
    .A2(_0265_),
    .B1(_0266_),
    .B2(_0267_),
    .X(_0268_));
 sky130_fd_sc_hd__or2_1 _1142_ (.A(net28),
    .B(net60),
    .X(_0269_));
 sky130_fd_sc_hd__nand2_1 _1143_ (.A(_0050_),
    .B(net60),
    .Y(_0270_));
 sky130_fd_sc_hd__xor2_2 _1144_ (.A(net26),
    .B(net58),
    .X(_0271_));
 sky130_fd_sc_hd__xor2_1 _1145_ (.A(net25),
    .B(net57),
    .X(_0272_));
 sky130_fd_sc_hd__xor2_4 _1146_ (.A(net61),
    .B(net29),
    .X(_0273_));
 sky130_fd_sc_hd__a2111oi_2 _1147_ (.A1(_0269_),
    .A2(_0270_),
    .B1(_0271_),
    .C1(_0272_),
    .D1(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__xnor2_1 _1148_ (.A(net22),
    .B(net54),
    .Y(_0275_));
 sky130_fd_sc_hd__or4bb_1 _1149_ (.A(_0263_),
    .B(_0268_),
    .C_N(_0274_),
    .D_N(_0275_),
    .X(_0276_));
 sky130_fd_sc_hd__buf_2 _1150_ (.A(net19),
    .X(_0277_));
 sky130_fd_sc_hd__nand2_1 _1151_ (.A(_0277_),
    .B(net51),
    .Y(_0278_));
 sky130_fd_sc_hd__or2_1 _1152_ (.A(net19),
    .B(net51),
    .X(_0279_));
 sky130_fd_sc_hd__xor2_1 _1153_ (.A(net20),
    .B(net52),
    .X(_0280_));
 sky130_fd_sc_hd__a21oi_1 _1154_ (.A1(_0278_),
    .A2(_0279_),
    .B1(_0280_),
    .Y(_0281_));
 sky130_fd_sc_hd__xnor2_1 _1155_ (.A(net18),
    .B(net50),
    .Y(_0282_));
 sky130_fd_sc_hd__xnor2_1 _1156_ (.A(net49),
    .B(net17),
    .Y(_0283_));
 sky130_fd_sc_hd__nand3_1 _1157_ (.A(_0281_),
    .B(_0282_),
    .C(_0283_),
    .Y(_0284_));
 sky130_fd_sc_hd__xor2_1 _1158_ (.A(net13),
    .B(net45),
    .X(_0285_));
 sky130_fd_sc_hd__or2_1 _1159_ (.A(net14),
    .B(net46),
    .X(_0286_));
 sky130_fd_sc_hd__buf_2 _1160_ (.A(net14),
    .X(_0287_));
 sky130_fd_sc_hd__nand2_1 _1161_ (.A(_0287_),
    .B(net46),
    .Y(_0288_));
 sky130_fd_sc_hd__buf_2 _1162_ (.A(net15),
    .X(_0289_));
 sky130_fd_sc_hd__xor2_1 _1163_ (.A(_0289_),
    .B(net47),
    .X(_0290_));
 sky130_fd_sc_hd__a21oi_1 _1164_ (.A1(_0286_),
    .A2(_0288_),
    .B1(_0290_),
    .Y(_0291_));
 sky130_fd_sc_hd__xnor2_1 _1165_ (.A(net44),
    .B(net12),
    .Y(_0292_));
 sky130_fd_sc_hd__nand2_1 _1166_ (.A(_0291_),
    .B(_0292_),
    .Y(_0293_));
 sky130_fd_sc_hd__or4_2 _1167_ (.A(_0276_),
    .B(_0284_),
    .C(_0285_),
    .D(_0293_),
    .X(_0294_));
 sky130_fd_sc_hd__a31o_1 _1168_ (.A1(_0242_),
    .A2(_0252_),
    .A3(_0260_),
    .B1(_0294_),
    .X(_0295_));
 sky130_fd_sc_hd__inv_2 _1169_ (.A(net13),
    .Y(_0296_));
 sky130_fd_sc_hd__buf_2 _1170_ (.A(net12),
    .X(_0297_));
 sky130_fd_sc_hd__nor2_1 _1171_ (.A(_0297_),
    .B(_0285_),
    .Y(_0298_));
 sky130_fd_sc_hd__a22o_1 _1172_ (.A1(_0296_),
    .A2(net45),
    .B1(net44),
    .B2(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__nand2_1 _1173_ (.A(_0291_),
    .B(_0299_),
    .Y(_0300_));
 sky130_fd_sc_hd__or3b_1 _1174_ (.A(_0287_),
    .B(_0290_),
    .C_N(net46),
    .X(_0301_));
 sky130_fd_sc_hd__inv_2 _1175_ (.A(_0289_),
    .Y(_0302_));
 sky130_fd_sc_hd__nand2_1 _1176_ (.A(_0302_),
    .B(net47),
    .Y(_0303_));
 sky130_fd_sc_hd__a31o_1 _1177_ (.A1(_0300_),
    .A2(_0301_),
    .A3(_0303_),
    .B1(_0284_),
    .X(_0304_));
 sky130_fd_sc_hd__or3b_1 _1178_ (.A(_0277_),
    .B(_0280_),
    .C_N(net51),
    .X(_0305_));
 sky130_fd_sc_hd__clkbuf_4 _1179_ (.A(net17),
    .X(_0306_));
 sky130_fd_sc_hd__inv_2 _1180_ (.A(_0306_),
    .Y(_0307_));
 sky130_fd_sc_hd__clkbuf_2 _1181_ (.A(net18),
    .X(_0308_));
 sky130_fd_sc_hd__and2b_1 _1182_ (.A_N(_0308_),
    .B(net50),
    .X(_0309_));
 sky130_fd_sc_hd__a31o_1 _1183_ (.A1(net49),
    .A2(_0307_),
    .A3(_0282_),
    .B1(_0309_),
    .X(_0310_));
 sky130_fd_sc_hd__clkbuf_2 _1184_ (.A(net20),
    .X(_0311_));
 sky130_fd_sc_hd__inv_2 _1185_ (.A(net52),
    .Y(_0312_));
 sky130_fd_sc_hd__o2bb2a_1 _1186_ (.A1_N(_0281_),
    .A2_N(_0310_),
    .B1(_0311_),
    .B2(_0312_),
    .X(_0313_));
 sky130_fd_sc_hd__a31o_1 _1187_ (.A1(_0304_),
    .A2(_0305_),
    .A3(_0313_),
    .B1(_0276_),
    .X(_0314_));
 sky130_fd_sc_hd__buf_2 _1188_ (.A(net24),
    .X(_0315_));
 sky130_fd_sc_hd__inv_2 _1189_ (.A(net56),
    .Y(_0316_));
 sky130_fd_sc_hd__buf_2 _1190_ (.A(net22),
    .X(_0317_));
 sky130_fd_sc_hd__inv_2 _1191_ (.A(_0317_),
    .Y(_0318_));
 sky130_fd_sc_hd__clkbuf_2 _1192_ (.A(net21),
    .X(_0319_));
 sky130_fd_sc_hd__and3b_1 _1193_ (.A_N(_0319_),
    .B(_0275_),
    .C(net53),
    .X(_0320_));
 sky130_fd_sc_hd__a21oi_1 _1194_ (.A1(_0318_),
    .A2(net54),
    .B1(_0320_),
    .Y(_0321_));
 sky130_fd_sc_hd__inv_2 _1195_ (.A(net55),
    .Y(_0322_));
 sky130_fd_sc_hd__a211o_1 _1196_ (.A1(_0264_),
    .A2(_0265_),
    .B1(_0119_),
    .C1(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__o221a_1 _1197_ (.A1(_0315_),
    .A2(_0316_),
    .B1(_0268_),
    .B2(_0321_),
    .C1(_0323_),
    .X(_0324_));
 sky130_fd_sc_hd__and2b_1 _1198_ (.A_N(_0324_),
    .B(_0274_),
    .X(_0325_));
 sky130_fd_sc_hd__inv_2 _1199_ (.A(_0325_),
    .Y(_0326_));
 sky130_fd_sc_hd__inv_2 _1200_ (.A(net61),
    .Y(_0327_));
 sky130_fd_sc_hd__buf_2 _1201_ (.A(net26),
    .X(_0328_));
 sky130_fd_sc_hd__or2b_1 _1202_ (.A(_0328_),
    .B_N(net58),
    .X(_0329_));
 sky130_fd_sc_hd__clkbuf_2 _1203_ (.A(net25),
    .X(_0330_));
 sky130_fd_sc_hd__or3b_1 _1204_ (.A(_0330_),
    .B(_0271_),
    .C_N(net57),
    .X(_0331_));
 sky130_fd_sc_hd__a221o_1 _1205_ (.A1(_0269_),
    .A2(_0270_),
    .B1(_0329_),
    .B2(_0331_),
    .C1(_0273_),
    .X(_0332_));
 sky130_fd_sc_hd__inv_2 _1206_ (.A(_0060_),
    .Y(_0333_));
 sky130_fd_sc_hd__clkbuf_4 _1207_ (.A(net1),
    .X(_0334_));
 sky130_fd_sc_hd__or4_1 _1208_ (.A(net61),
    .B(_0333_),
    .C(_0334_),
    .D(_0141_),
    .X(_0335_));
 sky130_fd_sc_hd__or3b_1 _1209_ (.A(_0050_),
    .B(_0273_),
    .C_N(net60),
    .X(_0336_));
 sky130_fd_sc_hd__o2111a_1 _1210_ (.A1(_0327_),
    .A2(_0060_),
    .B1(_0332_),
    .C1(_0335_),
    .D1(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__or2_1 _1211_ (.A(net16),
    .B(_0091_),
    .X(_0338_));
 sky130_fd_sc_hd__nand2_1 _1212_ (.A(_0159_),
    .B(_0091_),
    .Y(_0339_));
 sky130_fd_sc_hd__a2bb2o_1 _1213_ (.A1_N(_0180_),
    .A2_N(_0177_),
    .B1(_0338_),
    .B2(_0339_),
    .X(_0340_));
 sky130_fd_sc_hd__or3_1 _1214_ (.A(_0213_),
    .B(_0199_),
    .C(_0340_),
    .X(_0341_));
 sky130_fd_sc_hd__nor3_1 _1215_ (.A(_0294_),
    .B(_0241_),
    .C(_0341_),
    .Y(_0342_));
 sky130_fd_sc_hd__a31o_1 _1216_ (.A1(net61),
    .A2(_0333_),
    .A3(_0181_),
    .B1(_0141_),
    .X(_0343_));
 sky130_fd_sc_hd__or4b_1 _1217_ (.A(_0140_),
    .B(_0342_),
    .C(_0343_),
    .D_N(_0139_),
    .X(_0344_));
 sky130_fd_sc_hd__a41o_1 _1218_ (.A1(_0295_),
    .A2(_0314_),
    .A3(_0326_),
    .A4(_0337_),
    .B1(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__or2b_1 _1219_ (.A(_0191_),
    .B_N(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__clkbuf_1 _1220_ (.A(_0346_),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_4 _1221_ (.A(_0018_),
    .X(_0347_));
 sky130_fd_sc_hd__mux4_1 _1222_ (.A0(net18),
    .A1(_0277_),
    .A2(net20),
    .A3(_0319_),
    .S0(_0144_),
    .S1(_0193_),
    .X(_0348_));
 sky130_fd_sc_hd__mux4_1 _1223_ (.A0(net13),
    .A1(_0287_),
    .A2(_0289_),
    .A3(net17),
    .S0(_0144_),
    .S1(_0193_),
    .X(_0349_));
 sky130_fd_sc_hd__clkbuf_4 _1224_ (.A(_0125_),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _1225_ (.A0(_0348_),
    .A1(_0349_),
    .S(_0350_),
    .X(_0351_));
 sky130_fd_sc_hd__nor2_2 _1226_ (.A(_0135_),
    .B(_0170_),
    .Y(_0352_));
 sky130_fd_sc_hd__clkbuf_4 _1227_ (.A(_0124_),
    .X(_0353_));
 sky130_fd_sc_hd__mux4_1 _1228_ (.A0(_0317_),
    .A1(_0119_),
    .A2(_0315_),
    .A3(net25),
    .S0(_0144_),
    .S1(_0193_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _1229_ (.A0(_0328_),
    .A1(_0050_),
    .S(_0176_),
    .X(_0355_));
 sky130_fd_sc_hd__and2_1 _1230_ (.A(_0060_),
    .B(_0193_),
    .X(_0356_));
 sky130_fd_sc_hd__a21oi_1 _1231_ (.A1(_0160_),
    .A2(_0355_),
    .B1(_0356_),
    .Y(_0357_));
 sky130_fd_sc_hd__buf_4 _1232_ (.A(_0176_),
    .X(_0358_));
 sky130_fd_sc_hd__a21bo_1 _1233_ (.A1(_0050_),
    .A2(_0160_),
    .B1_N(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__nor2_1 _1234_ (.A(_0334_),
    .B(_0359_),
    .Y(_0360_));
 sky130_fd_sc_hd__o21ai_1 _1235_ (.A1(_0357_),
    .A2(_0360_),
    .B1(_0353_),
    .Y(_0361_));
 sky130_fd_sc_hd__o211a_1 _1236_ (.A1(_0353_),
    .A2(_0354_),
    .B1(_0361_),
    .C1(_0142_),
    .X(_0362_));
 sky130_fd_sc_hd__buf_2 _1237_ (.A(_0135_),
    .X(_0363_));
 sky130_fd_sc_hd__buf_2 _1238_ (.A(_0363_),
    .X(_0364_));
 sky130_fd_sc_hd__a22o_1 _1239_ (.A1(_0351_),
    .A2(_0352_),
    .B1(_0362_),
    .B2(_0364_),
    .X(_0365_));
 sky130_fd_sc_hd__or4b_1 _1240_ (.A(net2),
    .B(net3),
    .C(net4),
    .D_N(net1),
    .X(_0366_));
 sky130_fd_sc_hd__and3_1 _1241_ (.A(net48),
    .B(_0029_),
    .C(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__clkbuf_4 _1242_ (.A(_0366_),
    .X(_0368_));
 sky130_fd_sc_hd__a21oi_1 _1243_ (.A1(_0029_),
    .A2(_0368_),
    .B1(net48),
    .Y(_0369_));
 sky130_fd_sc_hd__or3_1 _1244_ (.A(net16),
    .B(_0367_),
    .C(_0369_),
    .X(_0370_));
 sky130_fd_sc_hd__o21ai_1 _1245_ (.A1(_0367_),
    .A2(_0369_),
    .B1(_0159_),
    .Y(_0371_));
 sky130_fd_sc_hd__nand2_1 _1246_ (.A(_0192_),
    .B(_0176_),
    .Y(_0372_));
 sky130_fd_sc_hd__a21oi_1 _1247_ (.A1(_0370_),
    .A2(_0371_),
    .B1(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__a311oi_1 _1248_ (.A1(_0370_),
    .A2(_0371_),
    .A3(_0372_),
    .B1(_0373_),
    .C1(_0185_),
    .Y(_0374_));
 sky130_fd_sc_hd__clkbuf_4 _1249_ (.A(_0154_),
    .X(_0375_));
 sky130_fd_sc_hd__clkbuf_4 _1250_ (.A(_0182_),
    .X(_0376_));
 sky130_fd_sc_hd__mux4_1 _1251_ (.A0(net9),
    .A1(net10),
    .A2(net11),
    .A3(net12),
    .S0(_0071_),
    .S1(_0091_),
    .X(_0377_));
 sky130_fd_sc_hd__mux4_1 _1252_ (.A0(net36),
    .A1(net6),
    .A2(net7),
    .A3(net8),
    .S0(_0071_),
    .S1(_0091_),
    .X(_0378_));
 sky130_fd_sc_hd__mux2_1 _1253_ (.A0(_0377_),
    .A1(_0378_),
    .S(_0125_),
    .X(_0379_));
 sky130_fd_sc_hd__mux4_1 _1254_ (.A0(_0159_),
    .A1(_0155_),
    .A2(_0156_),
    .A3(_0164_),
    .S0(_0144_),
    .S1(_0193_),
    .X(_0380_));
 sky130_fd_sc_hd__mux4_1 _1255_ (.A0(_0165_),
    .A1(_0166_),
    .A2(net34),
    .A3(_0232_),
    .S0(_0144_),
    .S1(_0193_),
    .X(_0381_));
 sky130_fd_sc_hd__nor2_1 _1256_ (.A(_0135_),
    .B(_0125_),
    .Y(_0382_));
 sky130_fd_sc_hd__a22o_1 _1257_ (.A1(_0152_),
    .A2(_0380_),
    .B1(_0381_),
    .B2(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__a21o_1 _1258_ (.A1(_0135_),
    .A2(_0379_),
    .B1(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__nor4b_1 _1259_ (.A(net1),
    .B(_0141_),
    .C(_0139_),
    .D_N(_0140_),
    .Y(_0385_));
 sky130_fd_sc_hd__and3_1 _1260_ (.A(net1),
    .B(_0141_),
    .C(_0178_),
    .X(_0386_));
 sky130_fd_sc_hd__buf_2 _1261_ (.A(_0386_),
    .X(_0387_));
 sky130_fd_sc_hd__a21o_1 _1262_ (.A1(_0385_),
    .A2(_0339_),
    .B1(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _1263_ (.A0(_0159_),
    .A1(net5),
    .S(_0144_),
    .X(_0389_));
 sky130_fd_sc_hd__nand2_1 _1264_ (.A(_0160_),
    .B(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__inv_2 _1265_ (.A(_0390_),
    .Y(_0391_));
 sky130_fd_sc_hd__and3_1 _1266_ (.A(_0174_),
    .B(_0152_),
    .C(_0391_),
    .X(_0392_));
 sky130_fd_sc_hd__a221o_1 _1267_ (.A1(_0171_),
    .A2(_0384_),
    .B1(_0388_),
    .B2(_0338_),
    .C1(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__a31o_1 _1268_ (.A1(_0159_),
    .A2(_0375_),
    .A3(_0376_),
    .B1(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__a211o_1 _1269_ (.A1(_0347_),
    .A2(_0365_),
    .B1(_0374_),
    .C1(_0394_),
    .X(net80));
 sky130_fd_sc_hd__and2b_1 _1270_ (.A_N(_0150_),
    .B(_0368_),
    .X(_0395_));
 sky130_fd_sc_hd__xnor2_1 _1271_ (.A(_0124_),
    .B(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__xnor2_1 _1272_ (.A(_0155_),
    .B(_0396_),
    .Y(_0397_));
 sky130_fd_sc_hd__a21boi_1 _1273_ (.A1(_0370_),
    .A2(_0372_),
    .B1_N(_0371_),
    .Y(_0398_));
 sky130_fd_sc_hd__nor2_1 _1274_ (.A(_0397_),
    .B(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hd__nand2_1 _1275_ (.A(_0397_),
    .B(_0398_),
    .Y(_0400_));
 sky130_fd_sc_hd__and2b_1 _1276_ (.A_N(_0141_),
    .B(_0178_),
    .X(_0401_));
 sky130_fd_sc_hd__clkbuf_4 _1277_ (.A(_0401_),
    .X(_0402_));
 sky130_fd_sc_hd__and3b_1 _1278_ (.A_N(_0399_),
    .B(_0400_),
    .C(_0402_),
    .X(_0403_));
 sky130_fd_sc_hd__mux2_1 _1279_ (.A0(_0155_),
    .A1(_0159_),
    .S(_0358_),
    .X(_0404_));
 sky130_fd_sc_hd__o21ai_2 _1280_ (.A1(_0375_),
    .A2(_0404_),
    .B1(_0194_),
    .Y(_0405_));
 sky130_fd_sc_hd__clkbuf_4 _1281_ (.A(_0385_),
    .X(_0406_));
 sky130_fd_sc_hd__a21oi_1 _1282_ (.A1(_0406_),
    .A2(_0198_),
    .B1(_0387_),
    .Y(_0407_));
 sky130_fd_sc_hd__nor2_1 _1283_ (.A(_0155_),
    .B(_0353_),
    .Y(_0408_));
 sky130_fd_sc_hd__mux2_1 _1284_ (.A0(net10),
    .A1(_0243_),
    .S(_0144_),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _1285_ (.A0(_0132_),
    .A1(_0409_),
    .S(_0160_),
    .X(_0410_));
 sky130_fd_sc_hd__mux4_1 _1286_ (.A0(_0253_),
    .A1(_0147_),
    .A2(_0248_),
    .A3(_0143_),
    .S0(_0157_),
    .S1(_0102_),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _1287_ (.A0(_0410_),
    .A1(_0411_),
    .S(_0350_),
    .X(_0412_));
 sky130_fd_sc_hd__mux4_1 _1288_ (.A0(_0155_),
    .A1(_0156_),
    .A2(_0164_),
    .A3(_0165_),
    .S0(_0157_),
    .S1(_0102_),
    .X(_0413_));
 sky130_fd_sc_hd__mux4_1 _1289_ (.A0(_0166_),
    .A1(_0167_),
    .A2(_0232_),
    .A3(_0146_),
    .S0(_0157_),
    .S1(_0102_),
    .X(_0414_));
 sky130_fd_sc_hd__a22o_1 _1290_ (.A1(_0152_),
    .A2(_0413_),
    .B1(_0414_),
    .B2(_0382_),
    .X(_0415_));
 sky130_fd_sc_hd__a21o_1 _1291_ (.A1(_0363_),
    .A2(_0412_),
    .B1(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__nand2_1 _1292_ (.A(_0171_),
    .B(_0416_),
    .Y(_0417_));
 sky130_fd_sc_hd__o221a_1 _1293_ (.A1(_0175_),
    .A2(_0405_),
    .B1(_0407_),
    .B2(_0408_),
    .C1(_0417_),
    .X(_0418_));
 sky130_fd_sc_hd__or4b_1 _1294_ (.A(net1),
    .B(_0140_),
    .C(_0139_),
    .D_N(_0141_),
    .X(_0419_));
 sky130_fd_sc_hd__clkbuf_4 _1295_ (.A(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__clkbuf_4 _1296_ (.A(_0137_),
    .X(_0421_));
 sky130_fd_sc_hd__nand2_1 _1297_ (.A(_0160_),
    .B(_0081_),
    .Y(_0422_));
 sky130_fd_sc_hd__nand2_1 _1298_ (.A(_0334_),
    .B(_0356_),
    .Y(_0423_));
 sky130_fd_sc_hd__mux2_1 _1299_ (.A0(_0039_),
    .A1(_0120_),
    .S(_0122_),
    .X(_0424_));
 sky130_fd_sc_hd__nor2_1 _1300_ (.A(_0353_),
    .B(_0424_),
    .Y(_0425_));
 sky130_fd_sc_hd__a31o_1 _1301_ (.A1(_0353_),
    .A2(_0422_),
    .A3(_0423_),
    .B1(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_1 _1302_ (.A0(_0121_),
    .A1(_0128_),
    .S(_0122_),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_1 _1303_ (.A0(_0129_),
    .A1(_0131_),
    .S(_0160_),
    .X(_0428_));
 sky130_fd_sc_hd__mux2_1 _1304_ (.A0(_0427_),
    .A1(_0428_),
    .S(_0350_),
    .X(_0429_));
 sky130_fd_sc_hd__nand2_1 _1305_ (.A(_0352_),
    .B(_0429_),
    .Y(_0430_));
 sky130_fd_sc_hd__o31a_1 _1306_ (.A1(_0421_),
    .A2(_0170_),
    .A3(_0426_),
    .B1(_0430_),
    .X(_0431_));
 sky130_fd_sc_hd__inv_2 _1307_ (.A(net63),
    .Y(_0432_));
 sky130_fd_sc_hd__o22a_1 _1308_ (.A1(_0420_),
    .A2(_0198_),
    .B1(_0431_),
    .B2(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__nand3b_1 _1309_ (.A_N(_0403_),
    .B(_0418_),
    .C(_0433_),
    .Y(net91));
 sky130_fd_sc_hd__and2_1 _1310_ (.A(_0155_),
    .B(_0396_),
    .X(_0434_));
 sky130_fd_sc_hd__o31a_1 _1311_ (.A1(net59),
    .A2(net48),
    .A3(_0029_),
    .B1(_0368_),
    .X(_0435_));
 sky130_fd_sc_hd__xnor2_1 _1312_ (.A(net62),
    .B(_0435_),
    .Y(_0436_));
 sky130_fd_sc_hd__xor2_2 _1313_ (.A(_0156_),
    .B(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__nand2_1 _1314_ (.A(_0434_),
    .B(_0437_),
    .Y(_0438_));
 sky130_fd_sc_hd__or3b_2 _1315_ (.A(_0397_),
    .B(_0398_),
    .C_N(_0437_),
    .X(_0439_));
 sky130_fd_sc_hd__and3_1 _1316_ (.A(_0402_),
    .B(_0438_),
    .C(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__o31a_1 _1317_ (.A1(_0434_),
    .A2(_0399_),
    .A3(_0437_),
    .B1(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__nor2_1 _1318_ (.A(_0181_),
    .B(_0170_),
    .Y(_0442_));
 sky130_fd_sc_hd__mux4_1 _1319_ (.A0(_0315_),
    .A1(_0330_),
    .A2(_0328_),
    .A3(_0050_),
    .S0(_0176_),
    .S1(_0193_),
    .X(_0443_));
 sky130_fd_sc_hd__and2_1 _1320_ (.A(_0126_),
    .B(_0443_),
    .X(_0444_));
 sky130_fd_sc_hd__nor2_1 _1321_ (.A(_0333_),
    .B(_0126_),
    .Y(_0445_));
 sky130_fd_sc_hd__or2_1 _1322_ (.A(_0444_),
    .B(_0445_),
    .X(_0446_));
 sky130_fd_sc_hd__mux4_1 _1323_ (.A0(_0311_),
    .A1(_0319_),
    .A2(_0317_),
    .A3(_0119_),
    .S0(_0176_),
    .S1(_0102_),
    .X(_0447_));
 sky130_fd_sc_hd__mux4_1 _1324_ (.A0(_0289_),
    .A1(net17),
    .A2(net18),
    .A3(_0277_),
    .S0(_0176_),
    .S1(_0193_),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _1325_ (.A0(_0447_),
    .A1(_0448_),
    .S(_0126_),
    .X(_0449_));
 sky130_fd_sc_hd__and2_1 _1326_ (.A(_0137_),
    .B(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__a21o_1 _1327_ (.A1(_0364_),
    .A2(_0446_),
    .B1(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__nor2_1 _1328_ (.A(_0334_),
    .B(_0170_),
    .Y(_0452_));
 sky130_fd_sc_hd__a31o_1 _1329_ (.A1(_0060_),
    .A2(_0353_),
    .A3(_0150_),
    .B1(_0444_),
    .X(_0453_));
 sky130_fd_sc_hd__a21o_1 _1330_ (.A1(_0364_),
    .A2(_0453_),
    .B1(_0450_),
    .X(_0454_));
 sky130_fd_sc_hd__a22o_1 _1331_ (.A1(_0442_),
    .A2(_0451_),
    .B1(_0452_),
    .B2(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__clkbuf_4 _1332_ (.A(_0171_),
    .X(_0456_));
 sky130_fd_sc_hd__mux4_1 _1333_ (.A0(_0243_),
    .A1(_0297_),
    .A2(net13),
    .A3(_0287_),
    .S0(_0358_),
    .S1(_0154_),
    .X(_0457_));
 sky130_fd_sc_hd__mux4_1 _1334_ (.A0(_0147_),
    .A1(_0248_),
    .A2(_0143_),
    .A3(_0245_),
    .S0(_0358_),
    .S1(_0154_),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _1335_ (.A0(_0457_),
    .A1(_0458_),
    .S(_0350_),
    .X(_0459_));
 sky130_fd_sc_hd__mux4_1 _1336_ (.A0(_0156_),
    .A1(_0164_),
    .A2(_0165_),
    .A3(_0166_),
    .S0(_0358_),
    .S1(_0154_),
    .X(_0460_));
 sky130_fd_sc_hd__mux4_1 _1337_ (.A0(_0167_),
    .A1(_0232_),
    .A2(_0146_),
    .A3(_0253_),
    .S0(_0358_),
    .S1(_0154_),
    .X(_0461_));
 sky130_fd_sc_hd__buf_2 _1338_ (.A(_0382_),
    .X(_0462_));
 sky130_fd_sc_hd__a22o_1 _1339_ (.A1(_0152_),
    .A2(_0460_),
    .B1(_0461_),
    .B2(_0462_),
    .X(_0463_));
 sky130_fd_sc_hd__a21o_1 _1340_ (.A1(_0364_),
    .A2(_0459_),
    .B1(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__mux4_2 _1341_ (.A0(_0156_),
    .A1(_0155_),
    .A2(_0159_),
    .A3(net5),
    .S0(_0176_),
    .S1(_0102_),
    .X(_0465_));
 sky130_fd_sc_hd__inv_2 _1342_ (.A(_0465_),
    .Y(_0466_));
 sky130_fd_sc_hd__nor2_1 _1343_ (.A(_0175_),
    .B(_0466_),
    .Y(_0467_));
 sky130_fd_sc_hd__and3_1 _1344_ (.A(_0385_),
    .B(_0195_),
    .C(_0196_),
    .X(_0468_));
 sky130_fd_sc_hd__a31o_1 _1345_ (.A1(_0156_),
    .A2(_0363_),
    .A3(_0376_),
    .B1(_0468_),
    .X(_0469_));
 sky130_fd_sc_hd__a211o_1 _1346_ (.A1(_0387_),
    .A2(_0195_),
    .B1(_0467_),
    .C1(_0469_),
    .X(_0470_));
 sky130_fd_sc_hd__a21o_1 _1347_ (.A1(_0456_),
    .A2(_0464_),
    .B1(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__a21oi_1 _1348_ (.A1(_0347_),
    .A2(_0455_),
    .B1(_0471_),
    .Y(_0472_));
 sky130_fd_sc_hd__or2b_1 _1349_ (.A(_0441_),
    .B_N(_0472_),
    .X(_0473_));
 sky130_fd_sc_hd__clkbuf_1 _1350_ (.A(_0473_),
    .X(net94));
 sky130_fd_sc_hd__and2_1 _1351_ (.A(_0156_),
    .B(_0436_),
    .X(_0474_));
 sky130_fd_sc_hd__a21oi_2 _1352_ (.A1(_0434_),
    .A2(_0437_),
    .B1(_0474_),
    .Y(_0475_));
 sky130_fd_sc_hd__or4_4 _1353_ (.A(net62),
    .B(net59),
    .C(net48),
    .D(net37),
    .X(_0476_));
 sky130_fd_sc_hd__nand2_1 _1354_ (.A(_0368_),
    .B(_0476_),
    .Y(_0477_));
 sky130_fd_sc_hd__xnor2_1 _1355_ (.A(_0432_),
    .B(_0477_),
    .Y(_0478_));
 sky130_fd_sc_hd__xnor2_1 _1356_ (.A(_0164_),
    .B(_0478_),
    .Y(_0479_));
 sky130_fd_sc_hd__a21oi_2 _1357_ (.A1(_0439_),
    .A2(_0475_),
    .B1(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__a31o_1 _1358_ (.A1(_0439_),
    .A2(_0475_),
    .A3(_0479_),
    .B1(_0185_),
    .X(_0481_));
 sky130_fd_sc_hd__a21o_1 _1359_ (.A1(_0350_),
    .A2(_0112_),
    .B1(_0445_),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _1360_ (.A0(_0123_),
    .A1(_0130_),
    .S(_0125_),
    .X(_0483_));
 sky130_fd_sc_hd__and2_1 _1361_ (.A(_0137_),
    .B(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__a21o_1 _1362_ (.A1(_0363_),
    .A2(_0482_),
    .B1(_0484_),
    .X(_0485_));
 sky130_fd_sc_hd__clkbuf_4 _1363_ (.A(_0126_),
    .X(_0486_));
 sky130_fd_sc_hd__a31o_1 _1364_ (.A1(_0363_),
    .A2(_0486_),
    .A3(_0112_),
    .B1(_0484_),
    .X(_0487_));
 sky130_fd_sc_hd__a22o_1 _1365_ (.A1(_0442_),
    .A2(_0485_),
    .B1(_0487_),
    .B2(_0452_),
    .X(_0488_));
 sky130_fd_sc_hd__clkbuf_4 _1366_ (.A(_0186_),
    .X(_0489_));
 sky130_fd_sc_hd__nand2_1 _1367_ (.A(_0136_),
    .B(_0174_),
    .Y(_0490_));
 sky130_fd_sc_hd__mux4_1 _1368_ (.A0(_0164_),
    .A1(net30),
    .A2(_0155_),
    .A3(_0159_),
    .S0(_0071_),
    .S1(_0091_),
    .X(_0491_));
 sky130_fd_sc_hd__nand2_1 _1369_ (.A(_0126_),
    .B(_0491_),
    .Y(_0492_));
 sky130_fd_sc_hd__o21ai_2 _1370_ (.A1(_0126_),
    .A2(_0151_),
    .B1(_0492_),
    .Y(_0493_));
 sky130_fd_sc_hd__or2b_1 _1371_ (.A(_0490_),
    .B_N(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__o221a_1 _1372_ (.A1(_0419_),
    .A2(_0210_),
    .B1(_0212_),
    .B2(_0489_),
    .C1(_0494_),
    .X(_0495_));
 sky130_fd_sc_hd__a21bo_1 _1373_ (.A1(_0387_),
    .A2(_0211_),
    .B1_N(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_1 _1374_ (.A0(_0133_),
    .A1(_0145_),
    .S(_0126_),
    .X(_0497_));
 sky130_fd_sc_hd__a22o_1 _1375_ (.A1(_0148_),
    .A2(_0382_),
    .B1(_0168_),
    .B2(_0152_),
    .X(_0498_));
 sky130_fd_sc_hd__a21o_1 _1376_ (.A1(_0363_),
    .A2(_0497_),
    .B1(_0498_),
    .X(_0499_));
 sky130_fd_sc_hd__and2_1 _1377_ (.A(_0171_),
    .B(_0499_),
    .X(_0500_));
 sky130_fd_sc_hd__a211o_1 _1378_ (.A1(_0347_),
    .A2(_0488_),
    .B1(_0496_),
    .C1(_0500_),
    .X(_0501_));
 sky130_fd_sc_hd__o21bai_1 _1379_ (.A1(_0480_),
    .A2(_0481_),
    .B1_N(_0501_),
    .Y(net95));
 sky130_fd_sc_hd__and2_1 _1380_ (.A(_0164_),
    .B(_0478_),
    .X(_0502_));
 sky130_fd_sc_hd__o21a_1 _1381_ (.A1(net63),
    .A2(_0476_),
    .B1(_0368_),
    .X(_0503_));
 sky130_fd_sc_hd__xnor2_2 _1382_ (.A(net64),
    .B(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__xnor2_1 _1383_ (.A(_0217_),
    .B(_0504_),
    .Y(_0505_));
 sky130_fd_sc_hd__o21ai_1 _1384_ (.A1(_0502_),
    .A2(_0480_),
    .B1(_0505_),
    .Y(_0506_));
 sky130_fd_sc_hd__or3_1 _1385_ (.A(_0502_),
    .B(_0480_),
    .C(_0505_),
    .X(_0507_));
 sky130_fd_sc_hd__nor2_1 _1386_ (.A(_0124_),
    .B(_0357_),
    .Y(_0508_));
 sky130_fd_sc_hd__or2_1 _1387_ (.A(_0445_),
    .B(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _1388_ (.A0(_0348_),
    .A1(_0354_),
    .S(_0124_),
    .X(_0510_));
 sky130_fd_sc_hd__and2_1 _1389_ (.A(_0137_),
    .B(_0510_),
    .X(_0511_));
 sky130_fd_sc_hd__a21o_1 _1390_ (.A1(_0363_),
    .A2(_0509_),
    .B1(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__a31o_1 _1391_ (.A1(_0363_),
    .A2(_0359_),
    .A3(_0508_),
    .B1(_0511_),
    .X(_0513_));
 sky130_fd_sc_hd__a22o_1 _1392_ (.A1(_0442_),
    .A2(_0512_),
    .B1(_0513_),
    .B2(_0452_),
    .X(_0514_));
 sky130_fd_sc_hd__clkbuf_4 _1393_ (.A(_0387_),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _1394_ (.A0(_0349_),
    .A1(_0377_),
    .S(_0126_),
    .X(_0516_));
 sky130_fd_sc_hd__and2_1 _1395_ (.A(_0152_),
    .B(_0381_),
    .X(_0517_));
 sky130_fd_sc_hd__a221o_1 _1396_ (.A1(_0382_),
    .A2(_0378_),
    .B1(_0516_),
    .B2(_0135_),
    .C1(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__and2_1 _1397_ (.A(_0171_),
    .B(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__mux2_1 _1398_ (.A0(net30),
    .A1(net27),
    .S(_0071_),
    .X(_0520_));
 sky130_fd_sc_hd__inv_2 _1399_ (.A(_0520_),
    .Y(_0521_));
 sky130_fd_sc_hd__mux2_1 _1400_ (.A0(_0217_),
    .A1(_0216_),
    .S(_0157_),
    .X(_0522_));
 sky130_fd_sc_hd__mux2_1 _1401_ (.A0(_0521_),
    .A1(_0522_),
    .S(_0160_),
    .X(_0523_));
 sky130_fd_sc_hd__mux2_2 _1402_ (.A0(_0390_),
    .A1(_0523_),
    .S(_0350_),
    .X(_0524_));
 sky130_fd_sc_hd__o22a_1 _1403_ (.A1(_0420_),
    .A2(_0207_),
    .B1(_0209_),
    .B2(_0489_),
    .X(_0525_));
 sky130_fd_sc_hd__o21ai_1 _1404_ (.A1(_0490_),
    .A2(_0524_),
    .B1(_0525_),
    .Y(_0526_));
 sky130_fd_sc_hd__a211o_1 _1405_ (.A1(_0515_),
    .A2(_0208_),
    .B1(_0519_),
    .C1(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__a21o_1 _1406_ (.A1(_0347_),
    .A2(_0514_),
    .B1(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__a31o_1 _1407_ (.A1(_0402_),
    .A2(_0506_),
    .A3(_0507_),
    .B1(_0528_),
    .X(net96));
 sky130_fd_sc_hd__o31a_1 _1408_ (.A1(net64),
    .A2(net63),
    .A3(_0476_),
    .B1(_0368_),
    .X(_0529_));
 sky130_fd_sc_hd__xnor2_1 _1409_ (.A(net65),
    .B(_0529_),
    .Y(_0530_));
 sky130_fd_sc_hd__xor2_1 _1410_ (.A(_0166_),
    .B(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__a21o_1 _1411_ (.A1(_0165_),
    .A2(_0504_),
    .B1(_0502_),
    .X(_0532_));
 sky130_fd_sc_hd__nor2_1 _1412_ (.A(_0165_),
    .B(_0504_),
    .Y(_0533_));
 sky130_fd_sc_hd__o21ba_1 _1413_ (.A1(_0480_),
    .A2(_0532_),
    .B1_N(_0533_),
    .X(_0534_));
 sky130_fd_sc_hd__nor2_1 _1414_ (.A(_0531_),
    .B(_0534_),
    .Y(_0535_));
 sky130_fd_sc_hd__o221a_1 _1415_ (.A1(_0165_),
    .A2(_0504_),
    .B1(_0532_),
    .B2(_0480_),
    .C1(_0531_),
    .X(_0536_));
 sky130_fd_sc_hd__a21o_1 _1416_ (.A1(_0406_),
    .A2(_0203_),
    .B1(_0515_),
    .X(_0537_));
 sky130_fd_sc_hd__nor2_1 _1417_ (.A(_0124_),
    .B(_0422_),
    .Y(_0538_));
 sky130_fd_sc_hd__or3_1 _1418_ (.A(_0356_),
    .B(_0445_),
    .C(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__mux2_1 _1419_ (.A0(_0427_),
    .A1(_0424_),
    .S(_0124_),
    .X(_0540_));
 sky130_fd_sc_hd__and2_1 _1420_ (.A(_0137_),
    .B(_0540_),
    .X(_0541_));
 sky130_fd_sc_hd__a21o_1 _1421_ (.A1(_0363_),
    .A2(_0539_),
    .B1(_0541_),
    .X(_0542_));
 sky130_fd_sc_hd__a21o_1 _1422_ (.A1(_0363_),
    .A2(_0538_),
    .B1(_0541_),
    .X(_0543_));
 sky130_fd_sc_hd__a22o_1 _1423_ (.A1(_0442_),
    .A2(_0542_),
    .B1(_0543_),
    .B2(_0452_),
    .X(_0544_));
 sky130_fd_sc_hd__mux2_1 _1424_ (.A0(_0428_),
    .A1(_0410_),
    .S(_0486_),
    .X(_0545_));
 sky130_fd_sc_hd__buf_2 _1425_ (.A(_0152_),
    .X(_0546_));
 sky130_fd_sc_hd__a22o_1 _1426_ (.A1(_0462_),
    .A2(_0411_),
    .B1(_0414_),
    .B2(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__a21o_1 _1427_ (.A1(_0364_),
    .A2(_0545_),
    .B1(_0547_),
    .X(_0548_));
 sky130_fd_sc_hd__mux4_1 _1428_ (.A0(_0166_),
    .A1(_0165_),
    .A2(_0164_),
    .A3(_0156_),
    .S0(_0157_),
    .S1(_0102_),
    .X(_0549_));
 sky130_fd_sc_hd__inv_2 _1429_ (.A(_0549_),
    .Y(_0550_));
 sky130_fd_sc_hd__mux2_1 _1430_ (.A0(_0405_),
    .A1(_0550_),
    .S(_0486_),
    .X(_0551_));
 sky130_fd_sc_hd__o22ai_1 _1431_ (.A1(_0420_),
    .A2(_0203_),
    .B1(_0551_),
    .B2(_0490_),
    .Y(_0552_));
 sky130_fd_sc_hd__a221o_1 _1432_ (.A1(_0347_),
    .A2(_0544_),
    .B1(_0548_),
    .B2(_0456_),
    .C1(_0552_),
    .X(_0553_));
 sky130_fd_sc_hd__a21oi_1 _1433_ (.A1(_0204_),
    .A2(_0537_),
    .B1(_0553_),
    .Y(_0554_));
 sky130_fd_sc_hd__o31ai_1 _1434_ (.A1(_0185_),
    .A2(_0535_),
    .A3(_0536_),
    .B1(_0554_),
    .Y(net97));
 sky130_fd_sc_hd__and2_1 _1435_ (.A(_0166_),
    .B(_0530_),
    .X(_0555_));
 sky130_fd_sc_hd__o41a_1 _1436_ (.A1(net65),
    .A2(net64),
    .A3(net63),
    .A4(_0476_),
    .B1(_0368_),
    .X(_0556_));
 sky130_fd_sc_hd__xnor2_2 _1437_ (.A(net66),
    .B(_0556_),
    .Y(_0557_));
 sky130_fd_sc_hd__xor2_1 _1438_ (.A(_0167_),
    .B(_0557_),
    .X(_0558_));
 sky130_fd_sc_hd__o21ai_1 _1439_ (.A1(_0555_),
    .A2(_0536_),
    .B1(_0558_),
    .Y(_0559_));
 sky130_fd_sc_hd__or3_1 _1440_ (.A(_0555_),
    .B(_0536_),
    .C(_0558_),
    .X(_0560_));
 sky130_fd_sc_hd__buf_2 _1441_ (.A(_0364_),
    .X(_0561_));
 sky130_fd_sc_hd__mux2_1 _1442_ (.A0(_0447_),
    .A1(_0443_),
    .S(_0353_),
    .X(_0562_));
 sky130_fd_sc_hd__and3_1 _1443_ (.A(_0060_),
    .B(_0486_),
    .C(_0150_),
    .X(_0563_));
 sky130_fd_sc_hd__nand2_1 _1444_ (.A(_0334_),
    .B(_0142_),
    .Y(_0564_));
 sky130_fd_sc_hd__nor2_2 _1445_ (.A(_0333_),
    .B(_0564_),
    .Y(_0565_));
 sky130_fd_sc_hd__a211o_1 _1446_ (.A1(_0452_),
    .A2(_0563_),
    .B1(_0565_),
    .C1(_0352_),
    .X(_0566_));
 sky130_fd_sc_hd__o21a_1 _1447_ (.A1(_0561_),
    .A2(_0562_),
    .B1(_0566_),
    .X(_0567_));
 sky130_fd_sc_hd__buf_2 _1448_ (.A(_0174_),
    .X(_0568_));
 sky130_fd_sc_hd__and2b_1 _1449_ (.A_N(_0176_),
    .B(net34),
    .X(_0569_));
 sky130_fd_sc_hd__a21oi_1 _1450_ (.A1(_0166_),
    .A2(_0358_),
    .B1(_0569_),
    .Y(_0570_));
 sky130_fd_sc_hd__mux2_1 _1451_ (.A0(_0522_),
    .A1(_0570_),
    .S(_0160_),
    .X(_0571_));
 sky130_fd_sc_hd__mux2_1 _1452_ (.A0(_0466_),
    .A1(_0571_),
    .S(_0486_),
    .X(_0572_));
 sky130_fd_sc_hd__inv_2 _1453_ (.A(_0572_),
    .Y(_0573_));
 sky130_fd_sc_hd__o21a_1 _1454_ (.A1(_0167_),
    .A2(net66),
    .B1(_0334_),
    .X(_0574_));
 sky130_fd_sc_hd__a21o_1 _1455_ (.A1(_0167_),
    .A2(net66),
    .B1(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__a32o_1 _1456_ (.A1(_0141_),
    .A2(_0178_),
    .A3(_0575_),
    .B1(_0205_),
    .B2(_0406_),
    .X(_0576_));
 sky130_fd_sc_hd__a31o_1 _1457_ (.A1(_0421_),
    .A2(_0568_),
    .A3(_0573_),
    .B1(_0576_),
    .X(_0577_));
 sky130_fd_sc_hd__mux2_1 _1458_ (.A0(_0448_),
    .A1(_0457_),
    .S(_0350_),
    .X(_0578_));
 sky130_fd_sc_hd__and2_1 _1459_ (.A(_0546_),
    .B(_0461_),
    .X(_0579_));
 sky130_fd_sc_hd__a221o_1 _1460_ (.A1(_0462_),
    .A2(_0458_),
    .B1(_0578_),
    .B2(_0364_),
    .C1(_0579_),
    .X(_0580_));
 sky130_fd_sc_hd__and2_1 _1461_ (.A(_0456_),
    .B(_0580_),
    .X(_0581_));
 sky130_fd_sc_hd__a211o_1 _1462_ (.A1(_0347_),
    .A2(_0567_),
    .B1(_0577_),
    .C1(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__a31o_1 _1463_ (.A1(_0402_),
    .A2(_0559_),
    .A3(_0560_),
    .B1(_0582_),
    .X(net98));
 sky130_fd_sc_hd__a22o_1 _1464_ (.A1(_0127_),
    .A2(_0352_),
    .B1(_0565_),
    .B2(_0364_),
    .X(_0583_));
 sky130_fd_sc_hd__mux2_1 _1465_ (.A0(_0134_),
    .A1(_0149_),
    .S(_0137_),
    .X(_0584_));
 sky130_fd_sc_hd__mux4_1 _1466_ (.A0(_0232_),
    .A1(net34),
    .A2(_0166_),
    .A3(_0165_),
    .S0(_0144_),
    .S1(_0193_),
    .X(_0585_));
 sky130_fd_sc_hd__mux2_1 _1467_ (.A0(_0491_),
    .A1(_0585_),
    .S(_0125_),
    .X(_0586_));
 sky130_fd_sc_hd__nand2_1 _1468_ (.A(_0135_),
    .B(_0126_),
    .Y(_0587_));
 sky130_fd_sc_hd__o2bb2a_1 _1469_ (.A1_N(_0137_),
    .A2_N(_0586_),
    .B1(_0587_),
    .B2(_0151_),
    .X(_0588_));
 sky130_fd_sc_hd__o2bb2a_1 _1470_ (.A1_N(_0142_),
    .A2_N(_0584_),
    .B1(_0588_),
    .B2(_0173_),
    .X(_0589_));
 sky130_fd_sc_hd__nor2_1 _1471_ (.A(_0018_),
    .B(_0589_),
    .Y(_0590_));
 sky130_fd_sc_hd__a221o_1 _1472_ (.A1(_0376_),
    .A2(_0231_),
    .B1(_0583_),
    .B2(_0018_),
    .C1(_0590_),
    .X(_0591_));
 sky130_fd_sc_hd__o21a_1 _1473_ (.A1(_0489_),
    .A2(_0231_),
    .B1(_0179_),
    .X(_0592_));
 sky130_fd_sc_hd__nor2_1 _1474_ (.A(_0233_),
    .B(_0592_),
    .Y(_0593_));
 sky130_fd_sc_hd__nand2_1 _1475_ (.A(_0531_),
    .B(_0558_),
    .Y(_0594_));
 sky130_fd_sc_hd__or2b_1 _1476_ (.A(_0479_),
    .B_N(_0505_),
    .X(_0595_));
 sky130_fd_sc_hd__a211o_1 _1477_ (.A1(_0439_),
    .A2(_0475_),
    .B1(_0594_),
    .C1(_0595_),
    .X(_0596_));
 sky130_fd_sc_hd__a21oi_1 _1478_ (.A1(_0165_),
    .A2(_0504_),
    .B1(_0502_),
    .Y(_0597_));
 sky130_fd_sc_hd__a21oi_1 _1479_ (.A1(_0167_),
    .A2(_0557_),
    .B1(_0555_),
    .Y(_0598_));
 sky130_fd_sc_hd__nor2_1 _1480_ (.A(_0167_),
    .B(_0557_),
    .Y(_0599_));
 sky130_fd_sc_hd__o32a_1 _1481_ (.A1(_0533_),
    .A2(_0597_),
    .A3(_0594_),
    .B1(_0598_),
    .B2(_0599_),
    .X(_0600_));
 sky130_fd_sc_hd__or4_2 _1482_ (.A(net66),
    .B(net65),
    .C(net64),
    .D(net63),
    .X(_0601_));
 sky130_fd_sc_hd__o21a_1 _1483_ (.A1(_0476_),
    .A2(_0601_),
    .B1(_0368_),
    .X(_0602_));
 sky130_fd_sc_hd__xnor2_1 _1484_ (.A(net67),
    .B(_0602_),
    .Y(_0603_));
 sky130_fd_sc_hd__and2_1 _1485_ (.A(_0232_),
    .B(_0603_),
    .X(_0604_));
 sky130_fd_sc_hd__nor2_1 _1486_ (.A(_0232_),
    .B(_0603_),
    .Y(_0605_));
 sky130_fd_sc_hd__or2_1 _1487_ (.A(_0604_),
    .B(_0605_),
    .X(_0606_));
 sky130_fd_sc_hd__and3_1 _1488_ (.A(_0596_),
    .B(_0600_),
    .C(_0606_),
    .X(_0607_));
 sky130_fd_sc_hd__a21oi_1 _1489_ (.A1(_0596_),
    .A2(_0600_),
    .B1(_0606_),
    .Y(_0608_));
 sky130_fd_sc_hd__or3_1 _1490_ (.A(_0185_),
    .B(_0607_),
    .C(_0608_),
    .X(_0609_));
 sky130_fd_sc_hd__or3b_1 _1491_ (.A(_0591_),
    .B(_0593_),
    .C_N(_0609_),
    .X(_0610_));
 sky130_fd_sc_hd__clkbuf_1 _1492_ (.A(_0610_),
    .X(net99));
 sky130_fd_sc_hd__buf_2 _1493_ (.A(_0368_),
    .X(_0611_));
 sky130_fd_sc_hd__clkbuf_4 _1494_ (.A(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__or3_1 _1495_ (.A(net67),
    .B(_0476_),
    .C(_0601_),
    .X(_0613_));
 sky130_fd_sc_hd__nand2_1 _1496_ (.A(_0612_),
    .B(_0613_),
    .Y(_0614_));
 sky130_fd_sc_hd__xor2_1 _1497_ (.A(net68),
    .B(_0614_),
    .X(_0615_));
 sky130_fd_sc_hd__xnor2_1 _1498_ (.A(_0255_),
    .B(_0615_),
    .Y(_0616_));
 sky130_fd_sc_hd__or3_1 _1499_ (.A(_0604_),
    .B(_0608_),
    .C(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__o21ai_1 _1500_ (.A1(_0604_),
    .A2(_0608_),
    .B1(_0616_),
    .Y(_0618_));
 sky130_fd_sc_hd__buf_2 _1501_ (.A(_0432_),
    .X(_0619_));
 sky130_fd_sc_hd__nand2_1 _1502_ (.A(_0364_),
    .B(_0565_),
    .Y(_0620_));
 sky130_fd_sc_hd__a21boi_1 _1503_ (.A1(_0421_),
    .A2(_0362_),
    .B1_N(_0620_),
    .Y(_0621_));
 sky130_fd_sc_hd__nor2_1 _1504_ (.A(_0619_),
    .B(_0621_),
    .Y(_0622_));
 sky130_fd_sc_hd__o21a_1 _1505_ (.A1(_0146_),
    .A2(net68),
    .B1(_0387_),
    .X(_0623_));
 sky130_fd_sc_hd__a31o_1 _1506_ (.A1(_0146_),
    .A2(net68),
    .A3(_0376_),
    .B1(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__and4bb_1 _1507_ (.A_N(_0141_),
    .B_N(_0139_),
    .C(_0140_),
    .D(net1),
    .X(_0625_));
 sky130_fd_sc_hd__buf_2 _1508_ (.A(_0625_),
    .X(_0626_));
 sky130_fd_sc_hd__nand2_2 _1509_ (.A(_0432_),
    .B(_0626_),
    .Y(_0627_));
 sky130_fd_sc_hd__inv_2 _1510_ (.A(net35),
    .Y(_0628_));
 sky130_fd_sc_hd__mux2_1 _1511_ (.A0(_0255_),
    .A1(_0628_),
    .S(_0157_),
    .X(_0629_));
 sky130_fd_sc_hd__mux2_1 _1512_ (.A0(_0570_),
    .A1(_0629_),
    .S(_0160_),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_1 _1513_ (.A0(_0523_),
    .A1(_0630_),
    .S(_0350_),
    .X(_0631_));
 sky130_fd_sc_hd__o22a_1 _1514_ (.A1(_0390_),
    .A2(_0587_),
    .B1(_0631_),
    .B2(_0364_),
    .X(_0632_));
 sky130_fd_sc_hd__mux2_1 _1515_ (.A0(_0351_),
    .A1(_0379_),
    .S(_0421_),
    .X(_0633_));
 sky130_fd_sc_hd__a2bb2o_1 _1516_ (.A1_N(_0627_),
    .A2_N(_0632_),
    .B1(_0633_),
    .B2(_0456_),
    .X(_0634_));
 sky130_fd_sc_hd__a2111o_1 _1517_ (.A1(_0406_),
    .A2(_0230_),
    .B1(_0622_),
    .C1(_0624_),
    .D1(_0634_),
    .X(_0635_));
 sky130_fd_sc_hd__a31o_1 _1518_ (.A1(_0402_),
    .A2(_0617_),
    .A3(_0618_),
    .B1(_0635_),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_4 _1519_ (.A(_0402_),
    .X(_0636_));
 sky130_fd_sc_hd__or4_2 _1520_ (.A(net68),
    .B(net67),
    .C(_0476_),
    .D(_0601_),
    .X(_0637_));
 sky130_fd_sc_hd__a21oi_1 _1521_ (.A1(_0612_),
    .A2(_0637_),
    .B1(net38),
    .Y(_0638_));
 sky130_fd_sc_hd__and3_1 _1522_ (.A(net38),
    .B(_0611_),
    .C(_0637_),
    .X(_0639_));
 sky130_fd_sc_hd__o21ai_1 _1523_ (.A1(_0638_),
    .A2(_0639_),
    .B1(_0253_),
    .Y(_0640_));
 sky130_fd_sc_hd__or3_1 _1524_ (.A(_0253_),
    .B(_0638_),
    .C(_0639_),
    .X(_0641_));
 sky130_fd_sc_hd__and2_1 _1525_ (.A(_0640_),
    .B(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__a21o_1 _1526_ (.A1(_0146_),
    .A2(_0615_),
    .B1(_0604_),
    .X(_0643_));
 sky130_fd_sc_hd__or2_1 _1527_ (.A(_0146_),
    .B(_0615_),
    .X(_0644_));
 sky130_fd_sc_hd__o21a_1 _1528_ (.A1(_0608_),
    .A2(_0643_),
    .B1(_0644_),
    .X(_0645_));
 sky130_fd_sc_hd__xor2_1 _1529_ (.A(_0642_),
    .B(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__and2_1 _1530_ (.A(_0387_),
    .B(_0235_),
    .X(_0647_));
 sky130_fd_sc_hd__a31o_1 _1531_ (.A1(_0406_),
    .A2(_0235_),
    .A3(_0236_),
    .B1(_0647_),
    .X(_0648_));
 sky130_fd_sc_hd__a31o_1 _1532_ (.A1(_0253_),
    .A2(net38),
    .A3(_0376_),
    .B1(_0648_),
    .X(_0649_));
 sky130_fd_sc_hd__clkbuf_4 _1533_ (.A(_0421_),
    .X(_0650_));
 sky130_fd_sc_hd__or2_1 _1534_ (.A(_0561_),
    .B(_0412_),
    .X(_0651_));
 sky130_fd_sc_hd__o211a_1 _1535_ (.A1(_0650_),
    .A2(_0429_),
    .B1(_0651_),
    .C1(_0456_),
    .X(_0652_));
 sky130_fd_sc_hd__clkbuf_4 _1536_ (.A(_0358_),
    .X(_0653_));
 sky130_fd_sc_hd__mux4_1 _1537_ (.A0(_0253_),
    .A1(_0146_),
    .A2(_0232_),
    .A3(_0167_),
    .S0(_0653_),
    .S1(_0375_),
    .X(_0654_));
 sky130_fd_sc_hd__mux2_1 _1538_ (.A0(_0549_),
    .A1(_0654_),
    .S(_0486_),
    .X(_0655_));
 sky130_fd_sc_hd__a2bb2o_1 _1539_ (.A1_N(_0405_),
    .A2_N(_0587_),
    .B1(_0655_),
    .B2(_0421_),
    .X(_0656_));
 sky130_fd_sc_hd__nand2_1 _1540_ (.A(_0421_),
    .B(_0142_),
    .Y(_0657_));
 sky130_fd_sc_hd__o21ai_1 _1541_ (.A1(_0657_),
    .A2(_0426_),
    .B1(_0620_),
    .Y(_0658_));
 sky130_fd_sc_hd__a22o_1 _1542_ (.A1(_0568_),
    .A2(_0656_),
    .B1(_0658_),
    .B2(_0347_),
    .X(_0659_));
 sky130_fd_sc_hd__or3_1 _1543_ (.A(_0649_),
    .B(_0652_),
    .C(_0659_),
    .X(_0660_));
 sky130_fd_sc_hd__a21o_1 _1544_ (.A1(_0636_),
    .A2(_0646_),
    .B1(_0660_),
    .X(net70));
 sky130_fd_sc_hd__o211ai_1 _1545_ (.A1(net38),
    .A2(_0637_),
    .B1(_0612_),
    .C1(_0258_),
    .Y(_0661_));
 sky130_fd_sc_hd__and2_1 _1546_ (.A(net38),
    .B(_0611_),
    .X(_0662_));
 sky130_fd_sc_hd__a211o_1 _1547_ (.A1(_0612_),
    .A2(_0637_),
    .B1(_0662_),
    .C1(_0258_),
    .X(_0663_));
 sky130_fd_sc_hd__nand3_1 _1548_ (.A(_0147_),
    .B(_0661_),
    .C(_0663_),
    .Y(_0664_));
 sky130_fd_sc_hd__a21o_1 _1549_ (.A1(_0661_),
    .A2(_0663_),
    .B1(_0147_),
    .X(_0665_));
 sky130_fd_sc_hd__and2_1 _1550_ (.A(_0664_),
    .B(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__a21boi_1 _1551_ (.A1(_0642_),
    .A2(_0645_),
    .B1_N(_0640_),
    .Y(_0667_));
 sky130_fd_sc_hd__xnor2_1 _1552_ (.A(_0666_),
    .B(_0667_),
    .Y(_0668_));
 sky130_fd_sc_hd__mux2_1 _1553_ (.A0(_0449_),
    .A1(_0459_),
    .S(_0650_),
    .X(_0669_));
 sky130_fd_sc_hd__clkbuf_4 _1554_ (.A(_0406_),
    .X(_0670_));
 sky130_fd_sc_hd__mux4_2 _1555_ (.A0(_0147_),
    .A1(_0253_),
    .A2(_0146_),
    .A3(_0232_),
    .S0(_0653_),
    .S1(_0154_),
    .X(_0671_));
 sky130_fd_sc_hd__inv_2 _1556_ (.A(_0671_),
    .Y(_0672_));
 sky130_fd_sc_hd__clkbuf_4 _1557_ (.A(_0486_),
    .X(_0673_));
 sky130_fd_sc_hd__mux2_1 _1558_ (.A0(_0571_),
    .A1(_0672_),
    .S(_0673_),
    .X(_0674_));
 sky130_fd_sc_hd__o22a_1 _1559_ (.A1(_0466_),
    .A2(_0587_),
    .B1(_0674_),
    .B2(_0561_),
    .X(_0675_));
 sky130_fd_sc_hd__nor2_1 _1560_ (.A(_0627_),
    .B(_0675_),
    .Y(_0676_));
 sky130_fd_sc_hd__clkbuf_4 _1561_ (.A(_0376_),
    .X(_0677_));
 sky130_fd_sc_hd__a2bb2o_1 _1562_ (.A1_N(_0179_),
    .A2_N(_0237_),
    .B1(_0238_),
    .B2(_0677_),
    .X(_0678_));
 sky130_fd_sc_hd__a211o_1 _1563_ (.A1(_0670_),
    .A2(_0239_),
    .B1(_0676_),
    .C1(_0678_),
    .X(_0679_));
 sky130_fd_sc_hd__buf_2 _1564_ (.A(_0561_),
    .X(_0680_));
 sky130_fd_sc_hd__nor2_1 _1565_ (.A(_0334_),
    .B(_0657_),
    .Y(_0681_));
 sky130_fd_sc_hd__a22o_1 _1566_ (.A1(_0680_),
    .A2(_0565_),
    .B1(_0681_),
    .B2(_0453_),
    .X(_0682_));
 sky130_fd_sc_hd__a31oi_2 _1567_ (.A1(_0334_),
    .A2(_0352_),
    .A3(_0446_),
    .B1(_0682_),
    .Y(_0683_));
 sky130_fd_sc_hd__nor2_1 _1568_ (.A(_0619_),
    .B(_0683_),
    .Y(_0684_));
 sky130_fd_sc_hd__a211o_1 _1569_ (.A1(_0456_),
    .A2(_0669_),
    .B1(_0679_),
    .C1(_0684_),
    .X(_0685_));
 sky130_fd_sc_hd__a21o_1 _1570_ (.A1(_0636_),
    .A2(_0668_),
    .B1(_0685_),
    .X(net71));
 sky130_fd_sc_hd__nand4b_1 _1571_ (.A_N(_0606_),
    .B(_0616_),
    .C(_0642_),
    .D(_0666_),
    .Y(_0686_));
 sky130_fd_sc_hd__a21o_1 _1572_ (.A1(_0596_),
    .A2(_0600_),
    .B1(_0686_),
    .X(_0687_));
 sky130_fd_sc_hd__a21boi_1 _1573_ (.A1(_0640_),
    .A2(_0664_),
    .B1_N(_0665_),
    .Y(_0688_));
 sky130_fd_sc_hd__a41o_1 _1574_ (.A1(_0644_),
    .A2(_0642_),
    .A3(_0643_),
    .A4(_0666_),
    .B1(_0688_),
    .X(_0689_));
 sky130_fd_sc_hd__inv_2 _1575_ (.A(_0689_),
    .Y(_0690_));
 sky130_fd_sc_hd__or4_1 _1576_ (.A(net39),
    .B(net38),
    .C(net68),
    .D(net67),
    .X(_0691_));
 sky130_fd_sc_hd__or3_1 _1577_ (.A(_0476_),
    .B(_0601_),
    .C(_0691_),
    .X(_0692_));
 sky130_fd_sc_hd__nand3b_1 _1578_ (.A_N(net40),
    .B(_0612_),
    .C(_0692_),
    .Y(_0693_));
 sky130_fd_sc_hd__a21bo_1 _1579_ (.A1(_0611_),
    .A2(_0692_),
    .B1_N(net40),
    .X(_0694_));
 sky130_fd_sc_hd__nand3_1 _1580_ (.A(_0248_),
    .B(_0693_),
    .C(_0694_),
    .Y(_0695_));
 sky130_fd_sc_hd__a21o_1 _1581_ (.A1(_0693_),
    .A2(_0694_),
    .B1(_0248_),
    .X(_0696_));
 sky130_fd_sc_hd__nand2_1 _1582_ (.A(_0695_),
    .B(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__a21o_1 _1583_ (.A1(_0687_),
    .A2(_0690_),
    .B1(_0697_),
    .X(_0698_));
 sky130_fd_sc_hd__nand3_1 _1584_ (.A(_0697_),
    .B(_0687_),
    .C(_0690_),
    .Y(_0699_));
 sky130_fd_sc_hd__a22oi_1 _1585_ (.A1(_0486_),
    .A2(_0112_),
    .B1(_0445_),
    .B2(_0334_),
    .Y(_0700_));
 sky130_fd_sc_hd__o21a_1 _1586_ (.A1(_0657_),
    .A2(_0700_),
    .B1(_0620_),
    .X(_0701_));
 sky130_fd_sc_hd__nor2_1 _1587_ (.A(_0432_),
    .B(_0701_),
    .Y(_0702_));
 sky130_fd_sc_hd__or2_1 _1588_ (.A(_0135_),
    .B(_0497_),
    .X(_0703_));
 sky130_fd_sc_hd__o211a_1 _1589_ (.A1(_0421_),
    .A2(_0483_),
    .B1(_0703_),
    .C1(_0171_),
    .X(_0704_));
 sky130_fd_sc_hd__a221o_1 _1590_ (.A1(_0515_),
    .A2(_0223_),
    .B1(_0225_),
    .B2(_0406_),
    .C1(_0704_),
    .X(_0705_));
 sky130_fd_sc_hd__mux4_1 _1591_ (.A0(_0248_),
    .A1(_0147_),
    .A2(_0253_),
    .A3(_0146_),
    .S0(_0157_),
    .S1(_0102_),
    .X(_0706_));
 sky130_fd_sc_hd__mux2_1 _1592_ (.A0(_0585_),
    .A1(_0706_),
    .S(_0350_),
    .X(_0707_));
 sky130_fd_sc_hd__mux2_1 _1593_ (.A0(_0493_),
    .A1(_0707_),
    .S(_0421_),
    .X(_0708_));
 sky130_fd_sc_hd__a2bb2o_1 _1594_ (.A1_N(_0420_),
    .A2_N(_0224_),
    .B1(_0708_),
    .B2(_0174_),
    .X(_0709_));
 sky130_fd_sc_hd__or3_1 _1595_ (.A(_0702_),
    .B(_0705_),
    .C(_0709_),
    .X(_0710_));
 sky130_fd_sc_hd__a31o_1 _1596_ (.A1(_0402_),
    .A2(_0698_),
    .A3(_0699_),
    .B1(_0710_),
    .X(net72));
 sky130_fd_sc_hd__or4_1 _1597_ (.A(net40),
    .B(_0476_),
    .C(_0601_),
    .D(_0691_),
    .X(_0711_));
 sky130_fd_sc_hd__clkbuf_2 _1598_ (.A(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__nand3_1 _1599_ (.A(net41),
    .B(_0612_),
    .C(_0712_),
    .Y(_0713_));
 sky130_fd_sc_hd__a21o_1 _1600_ (.A1(_0611_),
    .A2(_0712_),
    .B1(net41),
    .X(_0714_));
 sky130_fd_sc_hd__a21oi_1 _1601_ (.A1(_0713_),
    .A2(_0714_),
    .B1(_0247_),
    .Y(_0715_));
 sky130_fd_sc_hd__nand3_1 _1602_ (.A(_0247_),
    .B(_0713_),
    .C(_0714_),
    .Y(_0716_));
 sky130_fd_sc_hd__or2b_1 _1603_ (.A(_0715_),
    .B_N(_0716_),
    .X(_0717_));
 sky130_fd_sc_hd__nand3_1 _1604_ (.A(_0695_),
    .B(_0698_),
    .C(_0717_),
    .Y(_0718_));
 sky130_fd_sc_hd__a21o_1 _1605_ (.A1(_0695_),
    .A2(_0698_),
    .B1(_0717_),
    .X(_0719_));
 sky130_fd_sc_hd__and3_1 _1606_ (.A(_0636_),
    .B(_0718_),
    .C(_0719_),
    .X(_0720_));
 sky130_fd_sc_hd__mux2_1 _1607_ (.A0(_0516_),
    .A1(_0510_),
    .S(_0680_),
    .X(_0721_));
 sky130_fd_sc_hd__inv_2 _1608_ (.A(_0630_),
    .Y(_0722_));
 sky130_fd_sc_hd__mux4_1 _1609_ (.A0(_0143_),
    .A1(_0248_),
    .A2(_0147_),
    .A3(_0253_),
    .S0(_0653_),
    .S1(_0154_),
    .X(_0723_));
 sky130_fd_sc_hd__mux2_1 _1610_ (.A0(_0722_),
    .A1(_0723_),
    .S(_0486_),
    .X(_0724_));
 sky130_fd_sc_hd__nor2_1 _1611_ (.A(_0561_),
    .B(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hd__a211oi_1 _1612_ (.A1(_0680_),
    .A2(_0524_),
    .B1(_0725_),
    .C1(_0627_),
    .Y(_0726_));
 sky130_fd_sc_hd__o21a_1 _1613_ (.A1(_0143_),
    .A2(net41),
    .B1(_0515_),
    .X(_0727_));
 sky130_fd_sc_hd__a31o_1 _1614_ (.A1(_0143_),
    .A2(net41),
    .A3(_0376_),
    .B1(_0727_),
    .X(_0728_));
 sky130_fd_sc_hd__a211o_1 _1615_ (.A1(_0406_),
    .A2(_0222_),
    .B1(_0726_),
    .C1(_0728_),
    .X(_0729_));
 sky130_fd_sc_hd__and3_1 _1616_ (.A(_0359_),
    .B(_0508_),
    .C(_0681_),
    .X(_0730_));
 sky130_fd_sc_hd__a31o_1 _1617_ (.A1(_0334_),
    .A2(_0352_),
    .A3(_0509_),
    .B1(_0730_),
    .X(_0731_));
 sky130_fd_sc_hd__and2b_1 _1618_ (.A_N(_0731_),
    .B(_0620_),
    .X(_0732_));
 sky130_fd_sc_hd__nor2_1 _1619_ (.A(_0619_),
    .B(_0732_),
    .Y(_0733_));
 sky130_fd_sc_hd__a211o_1 _1620_ (.A1(_0456_),
    .A2(_0721_),
    .B1(_0729_),
    .C1(_0733_),
    .X(_0734_));
 sky130_fd_sc_hd__or2_1 _1621_ (.A(_0720_),
    .B(_0734_),
    .X(_0735_));
 sky130_fd_sc_hd__clkbuf_1 _1622_ (.A(_0735_),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_4 _1623_ (.A(_0185_),
    .X(_0736_));
 sky130_fd_sc_hd__o21a_1 _1624_ (.A1(net41),
    .A2(_0712_),
    .B1(_0611_),
    .X(_0737_));
 sky130_fd_sc_hd__xnor2_2 _1625_ (.A(net42),
    .B(_0737_),
    .Y(_0738_));
 sky130_fd_sc_hd__xor2_2 _1626_ (.A(_0245_),
    .B(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__inv_2 _1627_ (.A(_0739_),
    .Y(_0740_));
 sky130_fd_sc_hd__a41o_1 _1628_ (.A1(_0248_),
    .A2(_0693_),
    .A3(_0694_),
    .A4(_0716_),
    .B1(_0715_),
    .X(_0741_));
 sky130_fd_sc_hd__inv_2 _1629_ (.A(_0741_),
    .Y(_0742_));
 sky130_fd_sc_hd__or2_1 _1630_ (.A(_0698_),
    .B(_0717_),
    .X(_0743_));
 sky130_fd_sc_hd__and3_1 _1631_ (.A(_0740_),
    .B(_0742_),
    .C(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__a21oi_1 _1632_ (.A1(_0742_),
    .A2(_0743_),
    .B1(_0740_),
    .Y(_0745_));
 sky130_fd_sc_hd__o21a_1 _1633_ (.A1(_0245_),
    .A2(net42),
    .B1(_0515_),
    .X(_0746_));
 sky130_fd_sc_hd__a31o_1 _1634_ (.A1(_0245_),
    .A2(net42),
    .A3(_0677_),
    .B1(_0746_),
    .X(_0747_));
 sky130_fd_sc_hd__mux4_1 _1635_ (.A0(_0245_),
    .A1(_0143_),
    .A2(_0248_),
    .A3(_0147_),
    .S0(_0653_),
    .S1(_0375_),
    .X(_0748_));
 sky130_fd_sc_hd__or2_1 _1636_ (.A(_0673_),
    .B(_0654_),
    .X(_0749_));
 sky130_fd_sc_hd__o21ai_1 _1637_ (.A1(_0353_),
    .A2(_0748_),
    .B1(_0749_),
    .Y(_0750_));
 sky130_fd_sc_hd__mux2_1 _1638_ (.A0(_0551_),
    .A1(_0750_),
    .S(_0650_),
    .X(_0751_));
 sky130_fd_sc_hd__o22a_1 _1639_ (.A1(_0489_),
    .A2(_0227_),
    .B1(_0751_),
    .B2(_0627_),
    .X(_0752_));
 sky130_fd_sc_hd__mux2_1 _1640_ (.A0(_0540_),
    .A1(_0545_),
    .S(_0650_),
    .X(_0753_));
 sky130_fd_sc_hd__or2_1 _1641_ (.A(_0561_),
    .B(_0539_),
    .X(_0754_));
 sky130_fd_sc_hd__a21oi_1 _1642_ (.A1(_0333_),
    .A2(_0561_),
    .B1(_0564_),
    .Y(_0755_));
 sky130_fd_sc_hd__a22o_1 _1643_ (.A1(_0538_),
    .A2(_0681_),
    .B1(_0754_),
    .B2(_0755_),
    .X(_0756_));
 sky130_fd_sc_hd__clkbuf_4 _1644_ (.A(_0347_),
    .X(_0757_));
 sky130_fd_sc_hd__a22oi_2 _1645_ (.A1(_0456_),
    .A2(_0753_),
    .B1(_0756_),
    .B2(_0757_),
    .Y(_0758_));
 sky130_fd_sc_hd__and3b_1 _1646_ (.A_N(_0747_),
    .B(_0752_),
    .C(_0758_),
    .X(_0759_));
 sky130_fd_sc_hd__o31ai_1 _1647_ (.A1(_0736_),
    .A2(_0744_),
    .A3(_0745_),
    .B1(_0759_),
    .Y(net74));
 sky130_fd_sc_hd__and2_1 _1648_ (.A(_0245_),
    .B(_0738_),
    .X(_0760_));
 sky130_fd_sc_hd__o31a_1 _1649_ (.A1(net42),
    .A2(net41),
    .A3(_0712_),
    .B1(_0611_),
    .X(_0761_));
 sky130_fd_sc_hd__xnor2_1 _1650_ (.A(_0244_),
    .B(_0761_),
    .Y(_0762_));
 sky130_fd_sc_hd__xnor2_1 _1651_ (.A(_0243_),
    .B(_0762_),
    .Y(_0763_));
 sky130_fd_sc_hd__or3_1 _1652_ (.A(_0760_),
    .B(_0745_),
    .C(_0763_),
    .X(_0764_));
 sky130_fd_sc_hd__o21ai_1 _1653_ (.A1(_0760_),
    .A2(_0745_),
    .B1(_0763_),
    .Y(_0765_));
 sky130_fd_sc_hd__buf_2 _1654_ (.A(_0680_),
    .X(_0766_));
 sky130_fd_sc_hd__mux2_1 _1655_ (.A0(_0578_),
    .A1(_0562_),
    .S(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__and3_1 _1656_ (.A(_0243_),
    .B(net43),
    .C(_0677_),
    .X(_0768_));
 sky130_fd_sc_hd__inv_2 _1657_ (.A(_0243_),
    .Y(_0769_));
 sky130_fd_sc_hd__a21oi_1 _1658_ (.A1(_0769_),
    .A2(_0244_),
    .B1(_0179_),
    .Y(_0770_));
 sky130_fd_sc_hd__nand2_2 _1659_ (.A(_0347_),
    .B(_0565_),
    .Y(_0771_));
 sky130_fd_sc_hd__o21ai_1 _1660_ (.A1(_0489_),
    .A2(_0226_),
    .B1(_0771_),
    .Y(_0772_));
 sky130_fd_sc_hd__mux4_1 _1661_ (.A0(_0243_),
    .A1(_0245_),
    .A2(_0143_),
    .A3(_0248_),
    .S0(_0653_),
    .S1(_0375_),
    .X(_0773_));
 sky130_fd_sc_hd__mux2_1 _1662_ (.A0(_0671_),
    .A1(_0773_),
    .S(_0673_),
    .X(_0774_));
 sky130_fd_sc_hd__mux2_1 _1663_ (.A0(_0573_),
    .A1(_0774_),
    .S(_0650_),
    .X(_0775_));
 sky130_fd_sc_hd__a32o_1 _1664_ (.A1(_0757_),
    .A2(_0563_),
    .A3(_0681_),
    .B1(_0775_),
    .B2(_0568_),
    .X(_0776_));
 sky130_fd_sc_hd__or4_1 _1665_ (.A(_0768_),
    .B(_0770_),
    .C(_0772_),
    .D(_0776_),
    .X(_0777_));
 sky130_fd_sc_hd__a21o_1 _1666_ (.A1(_0456_),
    .A2(_0767_),
    .B1(_0777_),
    .X(_0778_));
 sky130_fd_sc_hd__a31o_1 _1667_ (.A1(_0636_),
    .A2(_0764_),
    .A3(_0765_),
    .B1(_0778_),
    .X(net75));
 sky130_fd_sc_hd__or4bb_1 _1668_ (.A(_0697_),
    .B(_0717_),
    .C_N(_0739_),
    .D_N(_0763_),
    .X(_0779_));
 sky130_fd_sc_hd__a211o_1 _1669_ (.A1(_0596_),
    .A2(_0600_),
    .B1(_0686_),
    .C1(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__and4bb_1 _1670_ (.A_N(_0697_),
    .B_N(_0717_),
    .C(_0739_),
    .D(_0763_),
    .X(_0781_));
 sky130_fd_sc_hd__a2bb2o_1 _1671_ (.A1_N(_0769_),
    .A2_N(_0762_),
    .B1(_0738_),
    .B2(_0245_),
    .X(_0782_));
 sky130_fd_sc_hd__nand2_1 _1672_ (.A(_0769_),
    .B(_0762_),
    .Y(_0783_));
 sky130_fd_sc_hd__a32o_1 _1673_ (.A1(_0739_),
    .A2(_0741_),
    .A3(_0763_),
    .B1(_0782_),
    .B2(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__a21oi_1 _1674_ (.A1(_0689_),
    .A2(_0781_),
    .B1(_0784_),
    .Y(_0785_));
 sky130_fd_sc_hd__or3_2 _1675_ (.A(net43),
    .B(net42),
    .C(net41),
    .X(_0786_));
 sky130_fd_sc_hd__o21a_1 _1676_ (.A1(_0712_),
    .A2(_0786_),
    .B1(_0611_),
    .X(_0787_));
 sky130_fd_sc_hd__xnor2_1 _1677_ (.A(net44),
    .B(_0787_),
    .Y(_0788_));
 sky130_fd_sc_hd__nand2_2 _1678_ (.A(_0297_),
    .B(_0788_),
    .Y(_0789_));
 sky130_fd_sc_hd__or2_1 _1679_ (.A(_0297_),
    .B(_0788_),
    .X(_0790_));
 sky130_fd_sc_hd__nand2_1 _1680_ (.A(_0789_),
    .B(_0790_),
    .Y(_0791_));
 sky130_fd_sc_hd__nand3_1 _1681_ (.A(_0780_),
    .B(_0785_),
    .C(_0791_),
    .Y(_0792_));
 sky130_fd_sc_hd__a21o_1 _1682_ (.A1(_0780_),
    .A2(_0785_),
    .B1(_0791_),
    .X(_0793_));
 sky130_fd_sc_hd__and3_1 _1683_ (.A(_0561_),
    .B(_0568_),
    .C(_0586_),
    .X(_0794_));
 sky130_fd_sc_hd__and3_1 _1684_ (.A(_0060_),
    .B(_0018_),
    .C(_0442_),
    .X(_0795_));
 sky130_fd_sc_hd__clkbuf_4 _1685_ (.A(_0795_),
    .X(_0796_));
 sky130_fd_sc_hd__a31o_1 _1686_ (.A1(net44),
    .A2(_0297_),
    .A3(_0376_),
    .B1(_0796_),
    .X(_0797_));
 sky130_fd_sc_hd__mux4_1 _1687_ (.A0(_0297_),
    .A1(_0243_),
    .A2(net10),
    .A3(_0143_),
    .S0(_0358_),
    .S1(_0154_),
    .X(_0798_));
 sky130_fd_sc_hd__mux2_1 _1688_ (.A0(_0706_),
    .A1(_0798_),
    .S(_0350_),
    .X(_0799_));
 sky130_fd_sc_hd__and3_1 _1689_ (.A(_0421_),
    .B(_0174_),
    .C(_0799_),
    .X(_0800_));
 sky130_fd_sc_hd__nor2_2 _1690_ (.A(_0432_),
    .B(_0173_),
    .Y(_0801_));
 sky130_fd_sc_hd__nand2_2 _1691_ (.A(_0137_),
    .B(_0801_),
    .Y(_0802_));
 sky130_fd_sc_hd__or2_1 _1692_ (.A(_0353_),
    .B(_0802_),
    .X(_0803_));
 sky130_fd_sc_hd__o21ai_1 _1693_ (.A1(net44),
    .A2(_0297_),
    .B1(_0387_),
    .Y(_0804_));
 sky130_fd_sc_hd__o221a_1 _1694_ (.A1(_0489_),
    .A2(_0292_),
    .B1(_0803_),
    .B2(_0151_),
    .C1(_0804_),
    .X(_0805_));
 sky130_fd_sc_hd__or3b_1 _1695_ (.A(_0797_),
    .B(_0800_),
    .C_N(_0805_),
    .X(_0806_));
 sky130_fd_sc_hd__a211o_1 _1696_ (.A1(_0138_),
    .A2(_0456_),
    .B1(_0794_),
    .C1(_0806_),
    .X(_0807_));
 sky130_fd_sc_hd__a31o_1 _1697_ (.A1(_0402_),
    .A2(_0792_),
    .A3(_0793_),
    .B1(_0807_),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_2 _1698_ (.A(net13),
    .X(_0808_));
 sky130_fd_sc_hd__o31a_1 _1699_ (.A1(net44),
    .A2(_0712_),
    .A3(_0786_),
    .B1(_0611_),
    .X(_0809_));
 sky130_fd_sc_hd__xnor2_1 _1700_ (.A(net45),
    .B(_0809_),
    .Y(_0810_));
 sky130_fd_sc_hd__nand2_1 _1701_ (.A(_0808_),
    .B(_0810_),
    .Y(_0811_));
 sky130_fd_sc_hd__or2_1 _1702_ (.A(_0808_),
    .B(_0810_),
    .X(_0812_));
 sky130_fd_sc_hd__nand2_1 _1703_ (.A(_0811_),
    .B(_0812_),
    .Y(_0813_));
 sky130_fd_sc_hd__nand3_1 _1704_ (.A(_0789_),
    .B(_0793_),
    .C(_0813_),
    .Y(_0814_));
 sky130_fd_sc_hd__a21o_1 _1705_ (.A1(_0789_),
    .A2(_0793_),
    .B1(_0813_),
    .X(_0815_));
 sky130_fd_sc_hd__inv_2 _1706_ (.A(_0802_),
    .Y(_0816_));
 sky130_fd_sc_hd__a21oi_1 _1707_ (.A1(_0808_),
    .A2(net45),
    .B1(_0489_),
    .Y(_0817_));
 sky130_fd_sc_hd__o22a_1 _1708_ (.A1(_0808_),
    .A2(net45),
    .B1(_0515_),
    .B2(_0817_),
    .X(_0818_));
 sky130_fd_sc_hd__a311o_1 _1709_ (.A1(_0808_),
    .A2(net45),
    .A3(_0376_),
    .B1(_0796_),
    .C1(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__mux4_1 _1710_ (.A0(_0808_),
    .A1(_0297_),
    .A2(_0243_),
    .A3(_0245_),
    .S0(_0358_),
    .S1(_0154_),
    .X(_0820_));
 sky130_fd_sc_hd__mux2_1 _1711_ (.A0(_0723_),
    .A1(_0820_),
    .S(_0486_),
    .X(_0821_));
 sky130_fd_sc_hd__nand2_1 _1712_ (.A(_0561_),
    .B(_0631_),
    .Y(_0822_));
 sky130_fd_sc_hd__o211a_1 _1713_ (.A1(_0561_),
    .A2(_0821_),
    .B1(_0822_),
    .C1(_0626_),
    .X(_0823_));
 sky130_fd_sc_hd__o21a_1 _1714_ (.A1(_0365_),
    .A2(_0823_),
    .B1(_0619_),
    .X(_0824_));
 sky130_fd_sc_hd__a311o_1 _1715_ (.A1(_0673_),
    .A2(_0391_),
    .A3(_0816_),
    .B1(_0819_),
    .C1(_0824_),
    .X(_0825_));
 sky130_fd_sc_hd__a31o_1 _1716_ (.A1(_0402_),
    .A2(_0814_),
    .A3(_0815_),
    .B1(_0825_),
    .X(net77));
 sky130_fd_sc_hd__nor2_1 _1717_ (.A(_0808_),
    .B(_0810_),
    .Y(_0826_));
 sky130_fd_sc_hd__and2_1 _1718_ (.A(net45),
    .B(_0368_),
    .X(_0827_));
 sky130_fd_sc_hd__or3_1 _1719_ (.A(net46),
    .B(_0809_),
    .C(_0827_),
    .X(_0828_));
 sky130_fd_sc_hd__o21ai_1 _1720_ (.A1(_0809_),
    .A2(_0827_),
    .B1(net46),
    .Y(_0829_));
 sky130_fd_sc_hd__inv_2 _1721_ (.A(_0287_),
    .Y(_0830_));
 sky130_fd_sc_hd__a21oi_1 _1722_ (.A1(_0828_),
    .A2(_0829_),
    .B1(_0830_),
    .Y(_0831_));
 sky130_fd_sc_hd__and3_1 _1723_ (.A(_0830_),
    .B(_0828_),
    .C(_0829_),
    .X(_0832_));
 sky130_fd_sc_hd__or2_1 _1724_ (.A(_0831_),
    .B(_0832_),
    .X(_0833_));
 sky130_fd_sc_hd__a311o_1 _1725_ (.A1(_0789_),
    .A2(_0793_),
    .A3(_0811_),
    .B1(_0826_),
    .C1(_0833_),
    .X(_0834_));
 sky130_fd_sc_hd__a31o_1 _1726_ (.A1(_0789_),
    .A2(_0793_),
    .A3(_0811_),
    .B1(_0826_),
    .X(_0835_));
 sky130_fd_sc_hd__a21oi_1 _1727_ (.A1(_0833_),
    .A2(_0835_),
    .B1(_0736_),
    .Y(_0836_));
 sky130_fd_sc_hd__a21oi_1 _1728_ (.A1(_0406_),
    .A2(_0288_),
    .B1(_0515_),
    .Y(_0837_));
 sky130_fd_sc_hd__nor2_1 _1729_ (.A(_0287_),
    .B(net46),
    .Y(_0838_));
 sky130_fd_sc_hd__o221a_1 _1730_ (.A1(_0420_),
    .A2(_0288_),
    .B1(_0837_),
    .B2(_0838_),
    .C1(_0771_),
    .X(_0839_));
 sky130_fd_sc_hd__mux4_1 _1731_ (.A0(_0287_),
    .A1(_0808_),
    .A2(_0297_),
    .A3(_0243_),
    .S0(_0653_),
    .S1(_0375_),
    .X(_0840_));
 sky130_fd_sc_hd__mux2_1 _1732_ (.A0(_0748_),
    .A1(_0840_),
    .S(_0673_),
    .X(_0841_));
 sky130_fd_sc_hd__o21a_1 _1733_ (.A1(_0650_),
    .A2(_0655_),
    .B1(_0626_),
    .X(_0842_));
 sky130_fd_sc_hd__o21ai_1 _1734_ (.A1(_0680_),
    .A2(_0841_),
    .B1(_0842_),
    .Y(_0843_));
 sky130_fd_sc_hd__a21o_1 _1735_ (.A1(_0431_),
    .A2(_0843_),
    .B1(_0347_),
    .X(_0844_));
 sky130_fd_sc_hd__o211a_1 _1736_ (.A1(_0405_),
    .A2(_0803_),
    .B1(_0839_),
    .C1(_0844_),
    .X(_0845_));
 sky130_fd_sc_hd__a21bo_1 _1737_ (.A1(_0834_),
    .A2(_0836_),
    .B1_N(_0845_),
    .X(_0846_));
 sky130_fd_sc_hd__clkbuf_1 _1738_ (.A(_0846_),
    .X(net78));
 sky130_fd_sc_hd__a21o_1 _1739_ (.A1(_0828_),
    .A2(_0829_),
    .B1(_0830_),
    .X(_0847_));
 sky130_fd_sc_hd__and2_1 _1740_ (.A(net46),
    .B(_0611_),
    .X(_0848_));
 sky130_fd_sc_hd__o31ai_1 _1741_ (.A1(_0809_),
    .A2(_0827_),
    .A3(_0848_),
    .B1(net47),
    .Y(_0849_));
 sky130_fd_sc_hd__a2111o_1 _1742_ (.A1(net46),
    .A2(_0612_),
    .B1(_0809_),
    .C1(_0827_),
    .D1(net47),
    .X(_0850_));
 sky130_fd_sc_hd__a21oi_1 _1743_ (.A1(_0849_),
    .A2(_0850_),
    .B1(_0302_),
    .Y(_0851_));
 sky130_fd_sc_hd__and3_1 _1744_ (.A(_0302_),
    .B(_0849_),
    .C(_0850_),
    .X(_0852_));
 sky130_fd_sc_hd__or2_1 _1745_ (.A(_0851_),
    .B(_0852_),
    .X(_0853_));
 sky130_fd_sc_hd__a21oi_1 _1746_ (.A1(_0847_),
    .A2(_0834_),
    .B1(_0853_),
    .Y(_0854_));
 sky130_fd_sc_hd__a31o_1 _1747_ (.A1(_0847_),
    .A2(_0834_),
    .A3(_0853_),
    .B1(_0736_),
    .X(_0855_));
 sky130_fd_sc_hd__nor2_1 _1748_ (.A(_0854_),
    .B(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__clkbuf_4 _1749_ (.A(_0653_),
    .X(_0857_));
 sky130_fd_sc_hd__buf_2 _1750_ (.A(_0375_),
    .X(_0858_));
 sky130_fd_sc_hd__mux4_1 _1751_ (.A0(_0289_),
    .A1(_0287_),
    .A2(_0808_),
    .A3(_0297_),
    .S0(_0857_),
    .S1(_0858_),
    .X(_0859_));
 sky130_fd_sc_hd__mux2_1 _1752_ (.A0(_0773_),
    .A1(_0859_),
    .S(_0673_),
    .X(_0860_));
 sky130_fd_sc_hd__nand2_1 _1753_ (.A(_0680_),
    .B(_0674_),
    .Y(_0861_));
 sky130_fd_sc_hd__o211a_1 _1754_ (.A1(_0766_),
    .A2(_0860_),
    .B1(_0861_),
    .C1(_0626_),
    .X(_0862_));
 sky130_fd_sc_hd__o21a_1 _1755_ (.A1(_0455_),
    .A2(_0862_),
    .B1(_0619_),
    .X(_0863_));
 sky130_fd_sc_hd__clkbuf_4 _1756_ (.A(_0515_),
    .X(_0864_));
 sky130_fd_sc_hd__o21a_1 _1757_ (.A1(_0289_),
    .A2(net47),
    .B1(_0864_),
    .X(_0865_));
 sky130_fd_sc_hd__a311o_1 _1758_ (.A1(_0289_),
    .A2(net47),
    .A3(_0677_),
    .B1(_0796_),
    .C1(_0865_),
    .X(_0866_));
 sky130_fd_sc_hd__a311o_1 _1759_ (.A1(_0546_),
    .A2(_0465_),
    .A3(_0801_),
    .B1(_0863_),
    .C1(_0866_),
    .X(_0867_));
 sky130_fd_sc_hd__a211o_1 _1760_ (.A1(_0670_),
    .A2(_0290_),
    .B1(_0856_),
    .C1(_0867_),
    .X(net79));
 sky130_fd_sc_hd__o21a_1 _1761_ (.A1(net49),
    .A2(_0306_),
    .B1(_0515_),
    .X(_0868_));
 sky130_fd_sc_hd__nor2_1 _1762_ (.A(_0489_),
    .B(_0283_),
    .Y(_0869_));
 sky130_fd_sc_hd__a311o_1 _1763_ (.A1(net49),
    .A2(_0306_),
    .A3(_0376_),
    .B1(_0868_),
    .C1(_0869_),
    .X(_0870_));
 sky130_fd_sc_hd__a211o_1 _1764_ (.A1(_0493_),
    .A2(_0816_),
    .B1(_0870_),
    .C1(_0796_),
    .X(_0871_));
 sky130_fd_sc_hd__mux4_1 _1765_ (.A0(_0306_),
    .A1(_0289_),
    .A2(_0287_),
    .A3(_0808_),
    .S0(_0653_),
    .S1(_0375_),
    .X(_0872_));
 sky130_fd_sc_hd__mux2_1 _1766_ (.A0(_0798_),
    .A1(_0872_),
    .S(_0673_),
    .X(_0873_));
 sky130_fd_sc_hd__mux2_1 _1767_ (.A0(_0707_),
    .A1(_0873_),
    .S(_0650_),
    .X(_0874_));
 sky130_fd_sc_hd__a21oi_1 _1768_ (.A1(_0626_),
    .A2(_0874_),
    .B1(_0488_),
    .Y(_0875_));
 sky130_fd_sc_hd__nor2_1 _1769_ (.A(_0757_),
    .B(_0875_),
    .Y(_0876_));
 sky130_fd_sc_hd__clkbuf_4 _1770_ (.A(_0612_),
    .X(_0877_));
 sky130_fd_sc_hd__or4_1 _1771_ (.A(net47),
    .B(net46),
    .C(net45),
    .D(net44),
    .X(_0878_));
 sky130_fd_sc_hd__or3_1 _1772_ (.A(_0712_),
    .B(_0786_),
    .C(_0878_),
    .X(_0879_));
 sky130_fd_sc_hd__nand2_1 _1773_ (.A(_0877_),
    .B(_0879_),
    .Y(_0880_));
 sky130_fd_sc_hd__xor2_2 _1774_ (.A(net49),
    .B(_0880_),
    .X(_0881_));
 sky130_fd_sc_hd__xnor2_2 _1775_ (.A(_0306_),
    .B(_0881_),
    .Y(_0882_));
 sky130_fd_sc_hd__a21o_1 _1776_ (.A1(_0789_),
    .A2(_0811_),
    .B1(_0826_),
    .X(_0883_));
 sky130_fd_sc_hd__nor2_1 _1777_ (.A(_0831_),
    .B(_0851_),
    .Y(_0884_));
 sky130_fd_sc_hd__o32a_1 _1778_ (.A1(_0833_),
    .A2(_0853_),
    .A3(_0883_),
    .B1(_0884_),
    .B2(_0852_),
    .X(_0885_));
 sky130_fd_sc_hd__or4_1 _1779_ (.A(_0791_),
    .B(_0813_),
    .C(_0833_),
    .D(_0853_),
    .X(_0886_));
 sky130_fd_sc_hd__a21o_1 _1780_ (.A1(_0780_),
    .A2(_0785_),
    .B1(_0886_),
    .X(_0887_));
 sky130_fd_sc_hd__a21oi_2 _1781_ (.A1(_0885_),
    .A2(_0887_),
    .B1(_0882_),
    .Y(_0888_));
 sky130_fd_sc_hd__a311o_1 _1782_ (.A1(_0882_),
    .A2(_0885_),
    .A3(_0887_),
    .B1(_0888_),
    .C1(_0185_),
    .X(_0889_));
 sky130_fd_sc_hd__or3b_1 _1783_ (.A(_0871_),
    .B(_0876_),
    .C_N(_0889_),
    .X(_0890_));
 sky130_fd_sc_hd__clkbuf_1 _1784_ (.A(_0890_),
    .X(net81));
 sky130_fd_sc_hd__o21a_1 _1785_ (.A1(net49),
    .A2(_0879_),
    .B1(_0612_),
    .X(_0891_));
 sky130_fd_sc_hd__xnor2_1 _1786_ (.A(net50),
    .B(_0891_),
    .Y(_0892_));
 sky130_fd_sc_hd__nand2_1 _1787_ (.A(_0308_),
    .B(_0892_),
    .Y(_0893_));
 sky130_fd_sc_hd__or2_1 _1788_ (.A(_0308_),
    .B(_0892_),
    .X(_0894_));
 sky130_fd_sc_hd__nand2_1 _1789_ (.A(_0893_),
    .B(_0894_),
    .Y(_0895_));
 sky130_fd_sc_hd__a21o_1 _1790_ (.A1(_0306_),
    .A2(_0881_),
    .B1(_0888_),
    .X(_0896_));
 sky130_fd_sc_hd__xnor2_1 _1791_ (.A(_0895_),
    .B(_0896_),
    .Y(_0897_));
 sky130_fd_sc_hd__o21a_1 _1792_ (.A1(_0308_),
    .A2(net50),
    .B1(_0864_),
    .X(_0898_));
 sky130_fd_sc_hd__a31o_1 _1793_ (.A1(_0308_),
    .A2(net50),
    .A3(_0677_),
    .B1(_0898_),
    .X(_0899_));
 sky130_fd_sc_hd__mux4_1 _1794_ (.A0(_0308_),
    .A1(_0306_),
    .A2(_0289_),
    .A3(_0287_),
    .S0(_0653_),
    .S1(_0375_),
    .X(_0900_));
 sky130_fd_sc_hd__mux2_1 _1795_ (.A0(_0820_),
    .A1(_0900_),
    .S(_0673_),
    .X(_0901_));
 sky130_fd_sc_hd__or2_1 _1796_ (.A(_0680_),
    .B(_0901_),
    .X(_0902_));
 sky130_fd_sc_hd__o211a_1 _1797_ (.A1(_0650_),
    .A2(_0724_),
    .B1(_0902_),
    .C1(_0626_),
    .X(_0903_));
 sky130_fd_sc_hd__o21a_1 _1798_ (.A1(_0514_),
    .A2(_0903_),
    .B1(_0619_),
    .X(_0904_));
 sky130_fd_sc_hd__o221a_1 _1799_ (.A1(_0489_),
    .A2(_0282_),
    .B1(_0524_),
    .B2(_0802_),
    .C1(_0771_),
    .X(_0905_));
 sky130_fd_sc_hd__or3b_1 _1800_ (.A(_0899_),
    .B(_0904_),
    .C_N(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__a21o_1 _1801_ (.A1(_0636_),
    .A2(_0897_),
    .B1(_0906_),
    .X(net82));
 sky130_fd_sc_hd__a22o_1 _1802_ (.A1(_0306_),
    .A2(_0881_),
    .B1(_0892_),
    .B2(_0308_),
    .X(_0907_));
 sky130_fd_sc_hd__or2_1 _1803_ (.A(net50),
    .B(net49),
    .X(_0908_));
 sky130_fd_sc_hd__or4_1 _1804_ (.A(_0712_),
    .B(_0786_),
    .C(_0878_),
    .D(_0908_),
    .X(_0909_));
 sky130_fd_sc_hd__nand2_1 _1805_ (.A(_0612_),
    .B(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__xor2_1 _1806_ (.A(net51),
    .B(_0910_),
    .X(_0911_));
 sky130_fd_sc_hd__xor2_1 _1807_ (.A(_0277_),
    .B(_0911_),
    .X(_0912_));
 sky130_fd_sc_hd__o211ai_2 _1808_ (.A1(_0888_),
    .A2(_0907_),
    .B1(_0912_),
    .C1(_0894_),
    .Y(_0913_));
 sky130_fd_sc_hd__o21a_1 _1809_ (.A1(_0888_),
    .A2(_0907_),
    .B1(_0894_),
    .X(_0914_));
 sky130_fd_sc_hd__or2_1 _1810_ (.A(_0912_),
    .B(_0914_),
    .X(_0915_));
 sky130_fd_sc_hd__mux4_1 _1811_ (.A0(_0277_),
    .A1(_0308_),
    .A2(_0306_),
    .A3(_0289_),
    .S0(_0857_),
    .S1(_0858_),
    .X(_0916_));
 sky130_fd_sc_hd__mux2_1 _1812_ (.A0(_0840_),
    .A1(_0916_),
    .S(_0673_),
    .X(_0917_));
 sky130_fd_sc_hd__nand2_1 _1813_ (.A(_0680_),
    .B(_0750_),
    .Y(_0918_));
 sky130_fd_sc_hd__o211a_1 _1814_ (.A1(_0766_),
    .A2(_0917_),
    .B1(_0918_),
    .C1(_0626_),
    .X(_0919_));
 sky130_fd_sc_hd__nor2_1 _1815_ (.A(_0544_),
    .B(_0919_),
    .Y(_0920_));
 sky130_fd_sc_hd__a21o_1 _1816_ (.A1(_0670_),
    .A2(_0278_),
    .B1(_0864_),
    .X(_0921_));
 sky130_fd_sc_hd__a21oi_1 _1817_ (.A1(_0279_),
    .A2(_0921_),
    .B1(_0796_),
    .Y(_0922_));
 sky130_fd_sc_hd__o221a_1 _1818_ (.A1(_0551_),
    .A2(_0802_),
    .B1(_0920_),
    .B2(_0757_),
    .C1(_0922_),
    .X(_0923_));
 sky130_fd_sc_hd__o21ai_1 _1819_ (.A1(_0420_),
    .A2(_0278_),
    .B1(_0923_),
    .Y(_0924_));
 sky130_fd_sc_hd__a31o_1 _1820_ (.A1(_0636_),
    .A2(_0913_),
    .A3(_0915_),
    .B1(_0924_),
    .X(net83));
 sky130_fd_sc_hd__nand2_1 _1821_ (.A(_0277_),
    .B(_0911_),
    .Y(_0925_));
 sky130_fd_sc_hd__o21a_1 _1822_ (.A1(net51),
    .A2(_0909_),
    .B1(_0877_),
    .X(_0926_));
 sky130_fd_sc_hd__xnor2_1 _1823_ (.A(net52),
    .B(_0926_),
    .Y(_0927_));
 sky130_fd_sc_hd__nor2_1 _1824_ (.A(_0311_),
    .B(_0927_),
    .Y(_0928_));
 sky130_fd_sc_hd__nand2_1 _1825_ (.A(_0311_),
    .B(_0927_),
    .Y(_0929_));
 sky130_fd_sc_hd__or2b_1 _1826_ (.A(_0928_),
    .B_N(_0929_),
    .X(_0930_));
 sky130_fd_sc_hd__a21oi_1 _1827_ (.A1(_0925_),
    .A2(_0913_),
    .B1(_0930_),
    .Y(_0931_));
 sky130_fd_sc_hd__a31o_1 _1828_ (.A1(_0925_),
    .A2(_0913_),
    .A3(_0930_),
    .B1(_0736_),
    .X(_0932_));
 sky130_fd_sc_hd__mux4_1 _1829_ (.A0(_0311_),
    .A1(_0277_),
    .A2(_0308_),
    .A3(_0306_),
    .S0(_0857_),
    .S1(_0858_),
    .X(_0933_));
 sky130_fd_sc_hd__mux2_1 _1830_ (.A0(_0859_),
    .A1(_0933_),
    .S(_0673_),
    .X(_0934_));
 sky130_fd_sc_hd__mux2_1 _1831_ (.A0(_0774_),
    .A1(_0934_),
    .S(_0650_),
    .X(_0935_));
 sky130_fd_sc_hd__a21oi_1 _1832_ (.A1(_0626_),
    .A2(_0935_),
    .B1(_0567_),
    .Y(_0936_));
 sky130_fd_sc_hd__or2_1 _1833_ (.A(_0311_),
    .B(net52),
    .X(_0937_));
 sky130_fd_sc_hd__a22o_1 _1834_ (.A1(_0864_),
    .A2(_0937_),
    .B1(_0280_),
    .B2(_0670_),
    .X(_0938_));
 sky130_fd_sc_hd__a311o_1 _1835_ (.A1(_0311_),
    .A2(net52),
    .A3(_0677_),
    .B1(_0796_),
    .C1(_0938_),
    .X(_0939_));
 sky130_fd_sc_hd__a21oi_1 _1836_ (.A1(_0573_),
    .A2(_0816_),
    .B1(_0939_),
    .Y(_0940_));
 sky130_fd_sc_hd__o21a_1 _1837_ (.A1(_0757_),
    .A2(_0936_),
    .B1(_0940_),
    .X(_0941_));
 sky130_fd_sc_hd__o21a_1 _1838_ (.A1(_0931_),
    .A2(_0932_),
    .B1(_0941_),
    .X(_0942_));
 sky130_fd_sc_hd__inv_2 _1839_ (.A(_0942_),
    .Y(net84));
 sky130_fd_sc_hd__inv_2 _1840_ (.A(net53),
    .Y(_0943_));
 sky130_fd_sc_hd__a21o_1 _1841_ (.A1(net52),
    .A2(_0877_),
    .B1(_0926_),
    .X(_0944_));
 sky130_fd_sc_hd__xnor2_1 _1842_ (.A(_0943_),
    .B(_0944_),
    .Y(_0945_));
 sky130_fd_sc_hd__and2b_1 _1843_ (.A_N(_0945_),
    .B(_0319_),
    .X(_0946_));
 sky130_fd_sc_hd__and2b_1 _1844_ (.A_N(_0319_),
    .B(_0945_),
    .X(_0947_));
 sky130_fd_sc_hd__nor2_1 _1845_ (.A(_0946_),
    .B(_0947_),
    .Y(_0948_));
 sky130_fd_sc_hd__and3b_1 _1846_ (.A_N(_0928_),
    .B(_0929_),
    .C(_0912_),
    .X(_0949_));
 sky130_fd_sc_hd__or3b_1 _1847_ (.A(_0882_),
    .B(_0895_),
    .C_N(_0949_),
    .X(_0950_));
 sky130_fd_sc_hd__or4b_1 _1848_ (.A(_0882_),
    .B(_0885_),
    .C(_0895_),
    .D_N(_0949_),
    .X(_0951_));
 sky130_fd_sc_hd__o21a_1 _1849_ (.A1(_0925_),
    .A2(_0928_),
    .B1(_0929_),
    .X(_0952_));
 sky130_fd_sc_hd__nand3_1 _1850_ (.A(_0894_),
    .B(_0907_),
    .C(_0949_),
    .Y(_0953_));
 sky130_fd_sc_hd__o2111a_2 _1851_ (.A1(_0887_),
    .A2(_0950_),
    .B1(_0951_),
    .C1(_0952_),
    .D1(_0953_),
    .X(_0954_));
 sky130_fd_sc_hd__and2b_1 _1852_ (.A_N(_0948_),
    .B(_0954_),
    .X(_0955_));
 sky130_fd_sc_hd__and2b_1 _1853_ (.A_N(_0954_),
    .B(_0948_),
    .X(_0956_));
 sky130_fd_sc_hd__mux4_1 _1854_ (.A0(_0319_),
    .A1(_0311_),
    .A2(_0277_),
    .A3(_0308_),
    .S0(_0653_),
    .S1(_0375_),
    .X(_0957_));
 sky130_fd_sc_hd__and2_1 _1855_ (.A(_0546_),
    .B(_0957_),
    .X(_0958_));
 sky130_fd_sc_hd__a221o_1 _1856_ (.A1(_0680_),
    .A2(_0799_),
    .B1(_0872_),
    .B2(_0462_),
    .C1(_0958_),
    .X(_0959_));
 sky130_fd_sc_hd__nand2_1 _1857_ (.A(_0757_),
    .B(_0626_),
    .Y(_0960_));
 sky130_fd_sc_hd__a2bb2o_1 _1858_ (.A1_N(_0588_),
    .A2_N(_0960_),
    .B1(_0583_),
    .B2(_0619_),
    .X(_0961_));
 sky130_fd_sc_hd__a22o_1 _1859_ (.A1(_0515_),
    .A2(_0261_),
    .B1(_0263_),
    .B2(_0406_),
    .X(_0962_));
 sky130_fd_sc_hd__a311o_1 _1860_ (.A1(net53),
    .A2(_0319_),
    .A3(_0677_),
    .B1(_0796_),
    .C1(_0962_),
    .X(_0963_));
 sky130_fd_sc_hd__a211oi_1 _1861_ (.A1(_0568_),
    .A2(_0959_),
    .B1(_0961_),
    .C1(_0963_),
    .Y(_0964_));
 sky130_fd_sc_hd__o31ai_2 _1862_ (.A1(_0736_),
    .A2(_0955_),
    .A3(_0956_),
    .B1(_0964_),
    .Y(net85));
 sky130_fd_sc_hd__inv_2 _1863_ (.A(net54),
    .Y(_0965_));
 sky130_fd_sc_hd__or4_1 _1864_ (.A(net53),
    .B(net52),
    .C(net51),
    .D(_0909_),
    .X(_0966_));
 sky130_fd_sc_hd__nand2_1 _1865_ (.A(_0877_),
    .B(_0966_),
    .Y(_0967_));
 sky130_fd_sc_hd__xnor2_1 _1866_ (.A(_0965_),
    .B(_0967_),
    .Y(_0968_));
 sky130_fd_sc_hd__and2_1 _1867_ (.A(_0317_),
    .B(_0968_),
    .X(_0969_));
 sky130_fd_sc_hd__or2_1 _1868_ (.A(_0317_),
    .B(_0968_),
    .X(_0970_));
 sky130_fd_sc_hd__and2b_1 _1869_ (.A_N(_0969_),
    .B(_0970_),
    .X(_0971_));
 sky130_fd_sc_hd__nor2_1 _1870_ (.A(_0946_),
    .B(_0956_),
    .Y(_0972_));
 sky130_fd_sc_hd__xnor2_1 _1871_ (.A(_0971_),
    .B(_0972_),
    .Y(_0973_));
 sky130_fd_sc_hd__mux4_1 _1872_ (.A0(_0317_),
    .A1(_0319_),
    .A2(_0311_),
    .A3(_0277_),
    .S0(_0857_),
    .S1(_0858_),
    .X(_0974_));
 sky130_fd_sc_hd__a22o_1 _1873_ (.A1(_0766_),
    .A2(_0821_),
    .B1(_0974_),
    .B2(_0546_),
    .X(_0975_));
 sky130_fd_sc_hd__a21oi_1 _1874_ (.A1(_0462_),
    .A2(_0900_),
    .B1(_0975_),
    .Y(_0976_));
 sky130_fd_sc_hd__nor2_1 _1875_ (.A(_0317_),
    .B(net54),
    .Y(_0977_));
 sky130_fd_sc_hd__o22a_1 _1876_ (.A1(_0179_),
    .A2(_0977_),
    .B1(_0275_),
    .B2(_0489_),
    .X(_0978_));
 sky130_fd_sc_hd__o311a_1 _1877_ (.A1(_0318_),
    .A2(_0965_),
    .A3(_0420_),
    .B1(_0771_),
    .C1(_0978_),
    .X(_0979_));
 sky130_fd_sc_hd__o221a_1 _1878_ (.A1(_0757_),
    .A2(_0621_),
    .B1(_0632_),
    .B2(_0960_),
    .C1(_0979_),
    .X(_0980_));
 sky130_fd_sc_hd__o21ai_1 _1879_ (.A1(_0627_),
    .A2(_0976_),
    .B1(_0980_),
    .Y(_0981_));
 sky130_fd_sc_hd__a21o_1 _1880_ (.A1(_0636_),
    .A2(_0973_),
    .B1(_0981_),
    .X(net86));
 sky130_fd_sc_hd__o21a_1 _1881_ (.A1(net54),
    .A2(_0966_),
    .B1(_0877_),
    .X(_0000_));
 sky130_fd_sc_hd__xnor2_1 _1882_ (.A(net55),
    .B(_0000_),
    .Y(_0001_));
 sky130_fd_sc_hd__xor2_1 _1883_ (.A(_0119_),
    .B(_0001_),
    .X(_0002_));
 sky130_fd_sc_hd__nand2_1 _1884_ (.A(_0948_),
    .B(_0971_),
    .Y(_0003_));
 sky130_fd_sc_hd__o21ai_1 _1885_ (.A1(_0946_),
    .A2(_0969_),
    .B1(_0970_),
    .Y(_0004_));
 sky130_fd_sc_hd__o21ai_1 _1886_ (.A1(_0954_),
    .A2(_0003_),
    .B1(_0004_),
    .Y(_0005_));
 sky130_fd_sc_hd__nand2_1 _1887_ (.A(_0002_),
    .B(_0005_),
    .Y(_0006_));
 sky130_fd_sc_hd__o21a_1 _1888_ (.A1(_0002_),
    .A2(_0005_),
    .B1(_0636_),
    .X(_0007_));
 sky130_fd_sc_hd__mux4_1 _1889_ (.A0(_0119_),
    .A1(_0317_),
    .A2(_0319_),
    .A3(_0311_),
    .S0(_0857_),
    .S1(_0858_),
    .X(_0008_));
 sky130_fd_sc_hd__and2_1 _1890_ (.A(_0546_),
    .B(_0008_),
    .X(_0009_));
 sky130_fd_sc_hd__a221o_1 _1891_ (.A1(_0680_),
    .A2(_0841_),
    .B1(_0916_),
    .B2(_0462_),
    .C1(_0009_),
    .X(_0010_));
 sky130_fd_sc_hd__a22o_1 _1892_ (.A1(_0656_),
    .A2(_0801_),
    .B1(_0010_),
    .B2(_0568_),
    .X(_0011_));
 sky130_fd_sc_hd__a21o_1 _1893_ (.A1(_0670_),
    .A2(_0267_),
    .B1(_0864_),
    .X(_0012_));
 sky130_fd_sc_hd__o2bb2a_1 _1894_ (.A1_N(_0266_),
    .A2_N(_0012_),
    .B1(_0267_),
    .B2(_0420_),
    .X(_0013_));
 sky130_fd_sc_hd__or3b_1 _1895_ (.A(_0011_),
    .B(_0796_),
    .C_N(_0013_),
    .X(_0014_));
 sky130_fd_sc_hd__and2_1 _1896_ (.A(_0619_),
    .B(_0658_),
    .X(_0015_));
 sky130_fd_sc_hd__a211o_1 _1897_ (.A1(_0006_),
    .A2(_0007_),
    .B1(_0014_),
    .C1(_0015_),
    .X(net87));
 sky130_fd_sc_hd__o31a_1 _1898_ (.A1(net55),
    .A2(net54),
    .A3(_0966_),
    .B1(_0877_),
    .X(_0016_));
 sky130_fd_sc_hd__xnor2_1 _1899_ (.A(_0316_),
    .B(_0016_),
    .Y(_0017_));
 sky130_fd_sc_hd__xnor2_1 _1900_ (.A(_0315_),
    .B(_0017_),
    .Y(_0019_));
 sky130_fd_sc_hd__nand2_1 _1901_ (.A(_0119_),
    .B(_0001_),
    .Y(_0020_));
 sky130_fd_sc_hd__a21bo_1 _1902_ (.A1(_0002_),
    .A2(_0005_),
    .B1_N(_0020_),
    .X(_0021_));
 sky130_fd_sc_hd__xnor2_1 _1903_ (.A(_0019_),
    .B(_0021_),
    .Y(_0022_));
 sky130_fd_sc_hd__a21o_1 _1904_ (.A1(_0670_),
    .A2(_0265_),
    .B1(_0864_),
    .X(_0023_));
 sky130_fd_sc_hd__o21ai_1 _1905_ (.A1(_0420_),
    .A2(_0265_),
    .B1(_0771_),
    .Y(_0024_));
 sky130_fd_sc_hd__a21oi_1 _1906_ (.A1(_0264_),
    .A2(_0023_),
    .B1(_0024_),
    .Y(_0025_));
 sky130_fd_sc_hd__mux4_1 _1907_ (.A0(_0315_),
    .A1(_0119_),
    .A2(_0317_),
    .A3(_0319_),
    .S0(_0857_),
    .S1(_0858_),
    .X(_0026_));
 sky130_fd_sc_hd__a22o_1 _1908_ (.A1(_0462_),
    .A2(_0933_),
    .B1(_0026_),
    .B2(_0546_),
    .X(_0027_));
 sky130_fd_sc_hd__a21oi_1 _1909_ (.A1(_0766_),
    .A2(_0860_),
    .B1(_0027_),
    .Y(_0028_));
 sky130_fd_sc_hd__o22a_1 _1910_ (.A1(_0675_),
    .A2(_0960_),
    .B1(_0028_),
    .B2(_0627_),
    .X(_0030_));
 sky130_fd_sc_hd__o211a_1 _1911_ (.A1(_0757_),
    .A2(_0683_),
    .B1(_0025_),
    .C1(_0030_),
    .X(_0031_));
 sky130_fd_sc_hd__o21ai_1 _1912_ (.A1(_0736_),
    .A2(_0022_),
    .B1(_0031_),
    .Y(net88));
 sky130_fd_sc_hd__o21a_1 _1913_ (.A1(net56),
    .A2(_0016_),
    .B1(_0877_),
    .X(_0032_));
 sky130_fd_sc_hd__xnor2_1 _1914_ (.A(net57),
    .B(_0032_),
    .Y(_0033_));
 sky130_fd_sc_hd__and2_1 _1915_ (.A(_0330_),
    .B(_0033_),
    .X(_0034_));
 sky130_fd_sc_hd__nor2_1 _1916_ (.A(_0330_),
    .B(_0033_),
    .Y(_0035_));
 sky130_fd_sc_hd__nor2_1 _1917_ (.A(_0034_),
    .B(_0035_),
    .Y(_0036_));
 sky130_fd_sc_hd__nand2_1 _1918_ (.A(_0002_),
    .B(_0019_),
    .Y(_0037_));
 sky130_fd_sc_hd__or2_1 _1919_ (.A(_0004_),
    .B(_0037_),
    .X(_0038_));
 sky130_fd_sc_hd__inv_2 _1920_ (.A(_0017_),
    .Y(_0040_));
 sky130_fd_sc_hd__a21bo_1 _1921_ (.A1(_0315_),
    .A2(_0040_),
    .B1_N(_0020_),
    .X(_0041_));
 sky130_fd_sc_hd__o21ai_1 _1922_ (.A1(_0315_),
    .A2(_0040_),
    .B1(_0041_),
    .Y(_0042_));
 sky130_fd_sc_hd__o311ai_4 _1923_ (.A1(_0954_),
    .A2(_0003_),
    .A3(_0037_),
    .B1(_0038_),
    .C1(_0042_),
    .Y(_0043_));
 sky130_fd_sc_hd__xnor2_1 _1924_ (.A(_0036_),
    .B(_0043_),
    .Y(_0044_));
 sky130_fd_sc_hd__mux4_1 _1925_ (.A0(_0330_),
    .A1(_0315_),
    .A2(_0119_),
    .A3(_0317_),
    .S0(_0857_),
    .S1(_0858_),
    .X(_0045_));
 sky130_fd_sc_hd__a22o_1 _1926_ (.A1(_0462_),
    .A2(_0957_),
    .B1(_0045_),
    .B2(_0546_),
    .X(_0046_));
 sky130_fd_sc_hd__or2_1 _1927_ (.A(_0330_),
    .B(net57),
    .X(_0047_));
 sky130_fd_sc_hd__a31o_1 _1928_ (.A1(_0330_),
    .A2(net57),
    .A3(_0677_),
    .B1(_0796_),
    .X(_0048_));
 sky130_fd_sc_hd__a221o_1 _1929_ (.A1(_0864_),
    .A2(_0047_),
    .B1(_0272_),
    .B2(_0670_),
    .C1(_0048_),
    .X(_0049_));
 sky130_fd_sc_hd__a31o_1 _1930_ (.A1(_0766_),
    .A2(_0568_),
    .A3(_0873_),
    .B1(_0049_),
    .X(_0051_));
 sky130_fd_sc_hd__a221o_1 _1931_ (.A1(_0708_),
    .A2(_0801_),
    .B1(_0046_),
    .B2(_0568_),
    .C1(_0051_),
    .X(_0052_));
 sky130_fd_sc_hd__o21ba_1 _1932_ (.A1(_0757_),
    .A2(_0701_),
    .B1_N(_0052_),
    .X(_0053_));
 sky130_fd_sc_hd__o21a_1 _1933_ (.A1(_0736_),
    .A2(_0044_),
    .B1(_0053_),
    .X(_0054_));
 sky130_fd_sc_hd__inv_2 _1934_ (.A(_0054_),
    .Y(net89));
 sky130_fd_sc_hd__a21oi_1 _1935_ (.A1(_0036_),
    .A2(_0043_),
    .B1(_0034_),
    .Y(_0055_));
 sky130_fd_sc_hd__o21a_1 _1936_ (.A1(net57),
    .A2(_0032_),
    .B1(_0877_),
    .X(_0056_));
 sky130_fd_sc_hd__xnor2_1 _1937_ (.A(net58),
    .B(_0056_),
    .Y(_0057_));
 sky130_fd_sc_hd__and2_1 _1938_ (.A(_0328_),
    .B(_0057_),
    .X(_0058_));
 sky130_fd_sc_hd__nor2_1 _1939_ (.A(_0328_),
    .B(_0057_),
    .Y(_0059_));
 sky130_fd_sc_hd__or2_1 _1940_ (.A(_0058_),
    .B(_0059_),
    .X(_0061_));
 sky130_fd_sc_hd__xnor2_1 _1941_ (.A(_0055_),
    .B(_0061_),
    .Y(_0062_));
 sky130_fd_sc_hd__a211o_1 _1942_ (.A1(_0766_),
    .A2(_0524_),
    .B1(_0725_),
    .C1(_0960_),
    .X(_0063_));
 sky130_fd_sc_hd__o21a_1 _1943_ (.A1(_0328_),
    .A2(net58),
    .B1(_0864_),
    .X(_0064_));
 sky130_fd_sc_hd__a31o_1 _1944_ (.A1(_0328_),
    .A2(net58),
    .A3(_0677_),
    .B1(_0796_),
    .X(_0065_));
 sky130_fd_sc_hd__mux4_1 _1945_ (.A0(_0328_),
    .A1(_0330_),
    .A2(_0315_),
    .A3(_0119_),
    .S0(_0857_),
    .S1(_0858_),
    .X(_0066_));
 sky130_fd_sc_hd__a22o_1 _1946_ (.A1(_0462_),
    .A2(_0974_),
    .B1(_0066_),
    .B2(_0546_),
    .X(_0067_));
 sky130_fd_sc_hd__a21oi_1 _1947_ (.A1(_0766_),
    .A2(_0901_),
    .B1(_0067_),
    .Y(_0068_));
 sky130_fd_sc_hd__nor2_1 _1948_ (.A(_0627_),
    .B(_0068_),
    .Y(_0069_));
 sky130_fd_sc_hd__a2111oi_1 _1949_ (.A1(_0670_),
    .A2(_0271_),
    .B1(_0064_),
    .C1(_0065_),
    .D1(_0069_),
    .Y(_0070_));
 sky130_fd_sc_hd__o211a_1 _1950_ (.A1(_0757_),
    .A2(_0732_),
    .B1(_0063_),
    .C1(_0070_),
    .X(_0072_));
 sky130_fd_sc_hd__o21ai_1 _1951_ (.A1(_0736_),
    .A2(_0062_),
    .B1(_0072_),
    .Y(net90));
 sky130_fd_sc_hd__a21o_1 _1952_ (.A1(net58),
    .A2(_0877_),
    .B1(_0056_),
    .X(_0073_));
 sky130_fd_sc_hd__xnor2_1 _1953_ (.A(net60),
    .B(_0073_),
    .Y(_0074_));
 sky130_fd_sc_hd__xor2_1 _1954_ (.A(_0050_),
    .B(_0074_),
    .X(_0075_));
 sky130_fd_sc_hd__inv_2 _1955_ (.A(_0059_),
    .Y(_0076_));
 sky130_fd_sc_hd__a211o_1 _1956_ (.A1(_0036_),
    .A2(_0043_),
    .B1(_0058_),
    .C1(_0034_),
    .X(_0077_));
 sky130_fd_sc_hd__and2_1 _1957_ (.A(_0076_),
    .B(_0077_),
    .X(_0078_));
 sky130_fd_sc_hd__xor2_1 _1958_ (.A(_0075_),
    .B(_0078_),
    .X(_0079_));
 sky130_fd_sc_hd__o21ai_1 _1959_ (.A1(_0420_),
    .A2(_0270_),
    .B1(_0771_),
    .Y(_0080_));
 sky130_fd_sc_hd__a21o_1 _1960_ (.A1(_0670_),
    .A2(_0270_),
    .B1(_0864_),
    .X(_0082_));
 sky130_fd_sc_hd__a2bb2o_1 _1961_ (.A1_N(_0751_),
    .A2_N(_0960_),
    .B1(_0082_),
    .B2(_0269_),
    .X(_0083_));
 sky130_fd_sc_hd__mux4_1 _1962_ (.A0(_0050_),
    .A1(_0328_),
    .A2(_0330_),
    .A3(_0315_),
    .S0(_0857_),
    .S1(_0858_),
    .X(_0084_));
 sky130_fd_sc_hd__and2_1 _1963_ (.A(_0546_),
    .B(_0084_),
    .X(_0085_));
 sky130_fd_sc_hd__a221o_1 _1964_ (.A1(_0766_),
    .A2(_0917_),
    .B1(_0008_),
    .B2(_0462_),
    .C1(_0085_),
    .X(_0086_));
 sky130_fd_sc_hd__a22oi_1 _1965_ (.A1(_0619_),
    .A2(_0756_),
    .B1(_0086_),
    .B2(_0568_),
    .Y(_0087_));
 sky130_fd_sc_hd__or3b_1 _1966_ (.A(_0080_),
    .B(_0083_),
    .C_N(_0087_),
    .X(_0088_));
 sky130_fd_sc_hd__a21o_1 _1967_ (.A1(_0636_),
    .A2(_0079_),
    .B1(_0088_),
    .X(net92));
 sky130_fd_sc_hd__a32o_1 _1968_ (.A1(_0076_),
    .A2(_0075_),
    .A3(_0077_),
    .B1(_0074_),
    .B2(_0050_),
    .X(_0089_));
 sky130_fd_sc_hd__o21a_1 _1969_ (.A1(net60),
    .A2(_0073_),
    .B1(_0877_),
    .X(_0090_));
 sky130_fd_sc_hd__xnor2_1 _1970_ (.A(_0273_),
    .B(_0090_),
    .Y(_0092_));
 sky130_fd_sc_hd__xnor2_1 _1971_ (.A(_0089_),
    .B(_0092_),
    .Y(_0093_));
 sky130_fd_sc_hd__nand2_1 _1972_ (.A(_0775_),
    .B(_0801_),
    .Y(_0094_));
 sky130_fd_sc_hd__or2_1 _1973_ (.A(_0650_),
    .B(_0934_),
    .X(_0095_));
 sky130_fd_sc_hd__mux4_1 _1974_ (.A0(_0060_),
    .A1(_0050_),
    .A2(_0328_),
    .A3(_0330_),
    .S0(_0857_),
    .S1(_0858_),
    .X(_0096_));
 sky130_fd_sc_hd__o31a_1 _1975_ (.A1(_0766_),
    .A2(_0353_),
    .A3(_0096_),
    .B1(_0568_),
    .X(_0097_));
 sky130_fd_sc_hd__o211a_1 _1976_ (.A1(_0163_),
    .A2(_0026_),
    .B1(_0095_),
    .C1(_0097_),
    .X(_0098_));
 sky130_fd_sc_hd__o22a_1 _1977_ (.A1(net61),
    .A2(_0060_),
    .B1(_0864_),
    .B2(_0565_),
    .X(_0099_));
 sky130_fd_sc_hd__and3_1 _1978_ (.A(net61),
    .B(_0060_),
    .C(_0677_),
    .X(_0100_));
 sky130_fd_sc_hd__and3_1 _1979_ (.A(_0619_),
    .B(_0563_),
    .C(_0681_),
    .X(_0101_));
 sky130_fd_sc_hd__a211o_1 _1980_ (.A1(_0670_),
    .A2(_0273_),
    .B1(_0100_),
    .C1(_0101_),
    .X(_0103_));
 sky130_fd_sc_hd__nor3_1 _1981_ (.A(_0098_),
    .B(_0099_),
    .C(_0103_),
    .Y(_0104_));
 sky130_fd_sc_hd__o211ai_1 _1982_ (.A1(_0736_),
    .A2(_0093_),
    .B1(_0094_),
    .C1(_0104_),
    .Y(net93));
 sky130_fd_sc_hd__nor4b_1 _1983_ (.A(net80),
    .B(net91),
    .C(_0441_),
    .D_N(_0472_),
    .Y(_0105_));
 sky130_fd_sc_hd__nor4b_1 _1984_ (.A(net69),
    .B(net95),
    .C(net96),
    .D_N(_0105_),
    .Y(_0106_));
 sky130_fd_sc_hd__or4b_1 _1985_ (.A(net97),
    .B(net98),
    .C(net99),
    .D_N(_0106_),
    .X(_0107_));
 sky130_fd_sc_hd__or2_1 _1986_ (.A(net70),
    .B(_0107_),
    .X(_0108_));
 sky130_fd_sc_hd__or3_1 _1987_ (.A(net100),
    .B(net72),
    .C(net76),
    .X(_0109_));
 sky130_fd_sc_hd__or4_1 _1988_ (.A(_0720_),
    .B(_0734_),
    .C(net77),
    .D(_0109_),
    .X(_0110_));
 sky130_fd_sc_hd__or4_1 _1989_ (.A(net71),
    .B(net81),
    .C(_0108_),
    .D(_0110_),
    .X(_0111_));
 sky130_fd_sc_hd__or3_1 _1990_ (.A(net74),
    .B(net78),
    .C(net85),
    .X(_0113_));
 sky130_fd_sc_hd__or4_1 _1991_ (.A(net75),
    .B(net82),
    .C(_0111_),
    .D(_0113_),
    .X(_0114_));
 sky130_fd_sc_hd__a211o_1 _1992_ (.A1(_0636_),
    .A2(_0973_),
    .B1(_0981_),
    .C1(net87),
    .X(_0115_));
 sky130_fd_sc_hd__or2_1 _1993_ (.A(net79),
    .B(net83),
    .X(_0116_));
 sky130_fd_sc_hd__o2111a_1 _1994_ (.A1(_0736_),
    .A2(_0022_),
    .B1(_0031_),
    .C1(_0054_),
    .D1(_0942_),
    .X(_0117_));
 sky130_fd_sc_hd__or4b_1 _1995_ (.A(_0114_),
    .B(_0115_),
    .C(_0116_),
    .D_N(_0117_),
    .X(_0118_));
 sky130_fd_sc_hd__nor4_1 _1996_ (.A(net90),
    .B(net92),
    .C(net93),
    .D(_0118_),
    .Y(net101));
 sky130_fd_sc_hd__conb_1 alu_103 (.LO(net103));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_359 ();
 sky130_fd_sc_hd__buf_2 input1 (.A(alu_op[0]),
    .X(net1));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(alu_op[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(alu_op[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(alu_op[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input5 (.A(op1[0]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(op1[10]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(op1[11]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(op1[12]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(op1[13]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(op1[14]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(op1[15]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(op1[16]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(op1[17]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(op1[18]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(op1[19]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(op1[1]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(op1[20]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(op1[21]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(op1[22]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(op1[23]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(op1[24]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(op1[25]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(op1[26]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(op1[27]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(op1[28]),
    .X(net25));
 sky130_fd_sc_hd__dlymetal6s2s_1 input26 (.A(op1[29]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(op1[2]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(op1[30]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(op1[31]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input30 (.A(op1[3]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(op1[4]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(op1[5]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(op1[6]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(op1[7]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(op1[8]),
    .X(net35));
 sky130_fd_sc_hd__dlymetal6s2s_1 input36 (.A(op1[9]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(op2[0]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(op2[10]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(op2[11]),
    .X(net39));
 sky130_fd_sc_hd__dlymetal6s2s_1 input40 (.A(op2[12]),
    .X(net40));
 sky130_fd_sc_hd__buf_2 input41 (.A(op2[13]),
    .X(net41));
 sky130_fd_sc_hd__buf_2 input42 (.A(op2[14]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(op2[15]),
    .X(net43));
 sky130_fd_sc_hd__buf_2 input44 (.A(op2[16]),
    .X(net44));
 sky130_fd_sc_hd__buf_2 input45 (.A(op2[17]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(op2[18]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(op2[19]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(op2[1]),
    .X(net48));
 sky130_fd_sc_hd__buf_2 input49 (.A(op2[20]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(op2[21]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(op2[22]),
    .X(net51));
 sky130_fd_sc_hd__buf_2 input52 (.A(op2[23]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(op2[24]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(op2[25]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(op2[26]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(op2[27]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 input57 (.A(op2[28]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(op2[29]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input59 (.A(op2[2]),
    .X(net59));
 sky130_fd_sc_hd__buf_1 input60 (.A(op2[30]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_4 input61 (.A(op2[31]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 input62 (.A(op2[3]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 input63 (.A(op2[4]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 input64 (.A(op2[5]),
    .X(net64));
 sky130_fd_sc_hd__dlymetal6s2s_1 input65 (.A(op2[6]),
    .X(net65));
 sky130_fd_sc_hd__buf_2 input66 (.A(op2[7]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 input67 (.A(op2[8]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 input68 (.A(op2[9]),
    .X(net68));
 sky130_fd_sc_hd__buf_1 output69 (.A(net69),
    .X(result[0]));
 sky130_fd_sc_hd__buf_1 output70 (.A(net70),
    .X(result[10]));
 sky130_fd_sc_hd__buf_1 output71 (.A(net71),
    .X(result[11]));
 sky130_fd_sc_hd__buf_1 output72 (.A(net72),
    .X(result[12]));
 sky130_fd_sc_hd__buf_1 output73 (.A(net73),
    .X(result[13]));
 sky130_fd_sc_hd__buf_1 output74 (.A(net74),
    .X(result[14]));
 sky130_fd_sc_hd__buf_1 output75 (.A(net75),
    .X(result[15]));
 sky130_fd_sc_hd__buf_1 output76 (.A(net76),
    .X(result[16]));
 sky130_fd_sc_hd__buf_1 output77 (.A(net77),
    .X(result[17]));
 sky130_fd_sc_hd__buf_1 output78 (.A(net78),
    .X(result[18]));
 sky130_fd_sc_hd__buf_1 output79 (.A(net79),
    .X(result[19]));
 sky130_fd_sc_hd__buf_1 output80 (.A(net80),
    .X(result[1]));
 sky130_fd_sc_hd__buf_1 output81 (.A(net81),
    .X(result[20]));
 sky130_fd_sc_hd__buf_1 output82 (.A(net82),
    .X(result[21]));
 sky130_fd_sc_hd__buf_1 output83 (.A(net83),
    .X(result[22]));
 sky130_fd_sc_hd__buf_1 output84 (.A(net84),
    .X(result[23]));
 sky130_fd_sc_hd__buf_1 output85 (.A(net85),
    .X(result[24]));
 sky130_fd_sc_hd__buf_1 output86 (.A(net86),
    .X(result[25]));
 sky130_fd_sc_hd__buf_1 output87 (.A(net87),
    .X(result[26]));
 sky130_fd_sc_hd__buf_1 output88 (.A(net88),
    .X(result[27]));
 sky130_fd_sc_hd__buf_1 output89 (.A(net89),
    .X(result[28]));
 sky130_fd_sc_hd__buf_1 output90 (.A(net90),
    .X(result[29]));
 sky130_fd_sc_hd__buf_1 output91 (.A(net91),
    .X(result[2]));
 sky130_fd_sc_hd__buf_1 output92 (.A(net92),
    .X(result[30]));
 sky130_fd_sc_hd__buf_1 output93 (.A(net93),
    .X(result[31]));
 sky130_fd_sc_hd__buf_1 output94 (.A(net94),
    .X(result[3]));
 sky130_fd_sc_hd__buf_1 output95 (.A(net95),
    .X(result[4]));
 sky130_fd_sc_hd__buf_1 output96 (.A(net96),
    .X(result[5]));
 sky130_fd_sc_hd__buf_1 output97 (.A(net97),
    .X(result[6]));
 sky130_fd_sc_hd__buf_1 output98 (.A(net98),
    .X(result[7]));
 sky130_fd_sc_hd__buf_1 output99 (.A(net99),
    .X(result[8]));
 sky130_fd_sc_hd__buf_1 output100 (.A(net100),
    .X(result[9]));
 sky130_fd_sc_hd__buf_1 output101 (.A(net101),
    .X(zero));
 sky130_fd_sc_hd__conb_1 alu_102 (.LO(net102));
 assign carry_out = net102;
 assign overflow = net103;
endmodule
